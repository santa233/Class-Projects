
module fft_8pt ( clk, reset_n, valid_in, valid_out, xi0_r, xi1_r, xi2_r, xi3_r, 
        xi4_r, xi5_r, xi6_r, xi7_r, xo0_r, xo1_r, xo2_r, xo3_r, xo4_r, xo5_r, 
        xo6_r, xo7_r, xi0_i, xi1_i, xi2_i, xi3_i, xi4_i, xi5_i, xi6_i, xi7_i, 
        xo0_i, xo1_i, xo2_i, xo3_i, xo4_i, xo5_i, xo6_i, xo7_i, W0_8_r, W1_8_r, 
        W2_8_r, W3_8_r, W0_8_i, W1_8_i, W2_8_i, W3_8_i );
  input [63:0] xi0_r;
  input [63:0] xi1_r;
  input [63:0] xi2_r;
  input [63:0] xi3_r;
  input [63:0] xi4_r;
  input [63:0] xi5_r;
  input [63:0] xi6_r;
  input [63:0] xi7_r;
  output [63:0] xo0_r;
  output [63:0] xo1_r;
  output [63:0] xo2_r;
  output [63:0] xo3_r;
  output [63:0] xo4_r;
  output [63:0] xo5_r;
  output [63:0] xo6_r;
  output [63:0] xo7_r;
  input [63:0] xi0_i;
  input [63:0] xi1_i;
  input [63:0] xi2_i;
  input [63:0] xi3_i;
  input [63:0] xi4_i;
  input [63:0] xi5_i;
  input [63:0] xi6_i;
  input [63:0] xi7_i;
  output [63:0] xo0_i;
  output [63:0] xo1_i;
  output [63:0] xo2_i;
  output [63:0] xo3_i;
  output [63:0] xo4_i;
  output [63:0] xo5_i;
  output [63:0] xo6_i;
  output [63:0] xo7_i;
  input [63:0] W0_8_r;
  input [63:0] W1_8_r;
  input [63:0] W2_8_r;
  input [63:0] W3_8_r;
  input [63:0] W0_8_i;
  input [63:0] W1_8_i;
  input [63:0] W2_8_i;
  input [63:0] W3_8_i;
  input clk, reset_n, valid_in;
  output valid_out;
  wire   valid_in_d1r, s2_3_tmp_i_0_, s2_7_tmp_i_0_, dp_cluster_0_N99,
         dp_cluster_0_N98, dp_cluster_0_N97, dp_cluster_0_N96,
         dp_cluster_0_N95, dp_cluster_0_N94, dp_cluster_0_N93,
         dp_cluster_0_N92, dp_cluster_0_N91, dp_cluster_0_N90,
         dp_cluster_0_N89, dp_cluster_0_N88, dp_cluster_0_N87,
         dp_cluster_0_N86, dp_cluster_0_N85, dp_cluster_0_N84,
         dp_cluster_0_N83, dp_cluster_0_N82, dp_cluster_0_N81,
         dp_cluster_0_N80, dp_cluster_0_N79, dp_cluster_0_N78,
         dp_cluster_0_N77, dp_cluster_0_N76, dp_cluster_0_N75,
         dp_cluster_0_N74, dp_cluster_0_N73, dp_cluster_0_N72,
         dp_cluster_0_N71, dp_cluster_0_N70, dp_cluster_0_N69,
         dp_cluster_0_N68, dp_cluster_0_N67, dp_cluster_0_N66,
         dp_cluster_0_N65, dp_cluster_0_N64, dp_cluster_0_N63,
         dp_cluster_0_N62, dp_cluster_0_N61, dp_cluster_0_N60,
         dp_cluster_0_N59, dp_cluster_0_N58, dp_cluster_0_N57,
         dp_cluster_0_N111, dp_cluster_0_N110, dp_cluster_0_N109,
         dp_cluster_0_N108, dp_cluster_0_N107, dp_cluster_0_N106,
         dp_cluster_0_N105, dp_cluster_0_N104, dp_cluster_0_N103,
         dp_cluster_0_N102, dp_cluster_0_N101, dp_cluster_0_N100,
         dp_cluster_1_N224, dp_cluster_1_N223, dp_cluster_1_N222,
         dp_cluster_1_N221, dp_cluster_1_N220, dp_cluster_1_N219,
         dp_cluster_1_N218, dp_cluster_1_N217, dp_cluster_1_N216,
         dp_cluster_1_N215, dp_cluster_1_N214, dp_cluster_1_N213,
         dp_cluster_1_N212, dp_cluster_1_N211, dp_cluster_1_N210,
         dp_cluster_1_N209, dp_cluster_1_N208, dp_cluster_1_N207,
         dp_cluster_1_N206, dp_cluster_1_N205, dp_cluster_1_N204,
         dp_cluster_1_N203, dp_cluster_1_N202, dp_cluster_1_N201,
         dp_cluster_1_N200, dp_cluster_1_N199, dp_cluster_1_N198,
         dp_cluster_1_N197, dp_cluster_1_N196, dp_cluster_1_N195,
         dp_cluster_1_N194, dp_cluster_1_N193, dp_cluster_1_N192,
         dp_cluster_1_N191, dp_cluster_1_N190, dp_cluster_1_N189,
         dp_cluster_1_N188, dp_cluster_1_N187, dp_cluster_1_N186,
         dp_cluster_1_N185, dp_cluster_1_N184, dp_cluster_1_N183,
         dp_cluster_1_N182, dp_cluster_1_N181, dp_cluster_1_N180,
         dp_cluster_1_N179, dp_cluster_1_N178, dp_cluster_1_N177,
         dp_cluster_1_N176, dp_cluster_1_N175, dp_cluster_1_N174,
         dp_cluster_1_N173, dp_cluster_1_N172, dp_cluster_1_N171,
         dp_cluster_1_N170, dp_cluster_1_N169, dp_cluster_2_N9,
         dp_cluster_2_N8, dp_cluster_2_N7, dp_cluster_2_N6, dp_cluster_2_N55,
         dp_cluster_2_N54, dp_cluster_2_N53, dp_cluster_2_N52,
         dp_cluster_2_N51, dp_cluster_2_N50, dp_cluster_2_N5, dp_cluster_2_N49,
         dp_cluster_2_N48, dp_cluster_2_N47, dp_cluster_2_N46,
         dp_cluster_2_N45, dp_cluster_2_N44, dp_cluster_2_N43,
         dp_cluster_2_N42, dp_cluster_2_N41, dp_cluster_2_N40, dp_cluster_2_N4,
         dp_cluster_2_N39, dp_cluster_2_N38, dp_cluster_2_N37,
         dp_cluster_2_N36, dp_cluster_2_N35, dp_cluster_2_N34,
         dp_cluster_2_N33, dp_cluster_2_N32, dp_cluster_2_N31,
         dp_cluster_2_N30, dp_cluster_2_N3, dp_cluster_2_N29, dp_cluster_2_N28,
         dp_cluster_2_N27, dp_cluster_2_N26, dp_cluster_2_N25,
         dp_cluster_2_N24, dp_cluster_2_N23, dp_cluster_2_N22,
         dp_cluster_2_N21, dp_cluster_2_N20, dp_cluster_2_N2, dp_cluster_2_N19,
         dp_cluster_2_N18, dp_cluster_2_N17, dp_cluster_2_N16,
         dp_cluster_2_N15, dp_cluster_2_N14, dp_cluster_2_N13,
         dp_cluster_2_N12, dp_cluster_2_N11, dp_cluster_2_N10, dp_cluster_2_N1,
         dp_cluster_3_N168, dp_cluster_3_N167, dp_cluster_3_N166,
         dp_cluster_3_N165, dp_cluster_3_N164, dp_cluster_3_N163,
         dp_cluster_3_N162, dp_cluster_3_N161, dp_cluster_3_N160,
         dp_cluster_3_N159, dp_cluster_3_N158, dp_cluster_3_N157,
         dp_cluster_3_N156, dp_cluster_3_N155, dp_cluster_3_N154,
         dp_cluster_3_N153, dp_cluster_3_N152, dp_cluster_3_N151,
         dp_cluster_3_N150, dp_cluster_3_N149, dp_cluster_3_N148,
         dp_cluster_3_N147, dp_cluster_3_N146, dp_cluster_3_N145,
         dp_cluster_3_N144, dp_cluster_3_N143, dp_cluster_3_N142,
         dp_cluster_3_N141, dp_cluster_3_N140, dp_cluster_3_N139,
         dp_cluster_3_N138, dp_cluster_3_N137, dp_cluster_3_N136,
         dp_cluster_3_N135, dp_cluster_3_N134, dp_cluster_3_N133,
         dp_cluster_3_N132, dp_cluster_3_N131, dp_cluster_3_N130,
         dp_cluster_3_N129, dp_cluster_3_N128, dp_cluster_3_N127,
         dp_cluster_3_N126, dp_cluster_3_N125, dp_cluster_3_N124,
         dp_cluster_3_N123, dp_cluster_3_N122, dp_cluster_3_N121,
         dp_cluster_3_N120, dp_cluster_3_N119, dp_cluster_3_N118,
         dp_cluster_3_N117, dp_cluster_3_N116, dp_cluster_3_N115,
         dp_cluster_3_N114, dp_cluster_3_N113, dp_cluster_3_mult_512_C415_n376,
         dp_cluster_3_mult_512_C415_n375, dp_cluster_3_mult_512_C415_n374,
         dp_cluster_3_mult_512_C415_n373, dp_cluster_3_mult_512_C415_n372,
         dp_cluster_3_mult_512_C415_n371, dp_cluster_3_mult_512_C415_n370,
         dp_cluster_3_mult_512_C415_n369, dp_cluster_3_mult_512_C415_n368,
         dp_cluster_3_mult_512_C415_n367, dp_cluster_3_mult_512_C415_n366,
         dp_cluster_3_mult_512_C415_n365, dp_cluster_3_mult_512_C415_n364,
         dp_cluster_3_mult_512_C415_n363, dp_cluster_3_mult_512_C415_n362,
         dp_cluster_3_mult_512_C415_n361, dp_cluster_3_mult_512_C415_n360,
         dp_cluster_3_mult_512_C415_n359, dp_cluster_3_mult_512_C415_n358,
         dp_cluster_3_mult_512_C415_n357, dp_cluster_3_mult_512_C415_n356,
         dp_cluster_3_mult_512_C415_n355, dp_cluster_3_mult_512_C415_n354,
         dp_cluster_3_mult_512_C415_n353, dp_cluster_3_mult_512_C415_n352,
         dp_cluster_3_mult_512_C415_n351, dp_cluster_3_mult_512_C415_n350,
         dp_cluster_3_mult_512_C415_n349, dp_cluster_3_mult_512_C415_n348,
         dp_cluster_3_mult_512_C415_n347, dp_cluster_3_mult_512_C415_n346,
         dp_cluster_3_mult_512_C415_n345, dp_cluster_3_mult_512_C415_n344,
         dp_cluster_3_mult_512_C415_n343, dp_cluster_3_mult_512_C415_n342,
         dp_cluster_3_mult_512_C415_n341, dp_cluster_3_mult_512_C415_n340,
         dp_cluster_3_mult_512_C415_n339, dp_cluster_3_mult_512_C415_n338,
         dp_cluster_3_mult_512_C415_n337, dp_cluster_3_mult_512_C415_n336,
         dp_cluster_3_mult_512_C415_n335, dp_cluster_3_mult_512_C415_n334,
         dp_cluster_3_mult_512_C415_n333, dp_cluster_3_mult_512_C415_n332,
         dp_cluster_3_mult_512_C415_n331, dp_cluster_3_mult_512_C415_n330,
         dp_cluster_3_mult_512_C415_n329, dp_cluster_3_mult_512_C415_n328,
         dp_cluster_3_mult_512_C415_n327, dp_cluster_3_mult_512_C415_n326,
         dp_cluster_3_mult_512_C415_n325, dp_cluster_3_mult_512_C415_n324,
         dp_cluster_3_mult_512_C415_n323, dp_cluster_3_mult_512_C415_n322,
         dp_cluster_3_mult_512_C415_n321, dp_cluster_3_mult_512_C415_n320,
         dp_cluster_3_mult_512_C415_n319, dp_cluster_3_mult_512_C415_n317,
         dp_cluster_3_mult_512_C415_n316, dp_cluster_3_mult_512_C415_n315,
         dp_cluster_3_mult_512_C415_n314, dp_cluster_3_mult_512_C415_n313,
         dp_cluster_3_mult_512_C415_n312, dp_cluster_3_mult_512_C415_n311,
         dp_cluster_3_mult_512_C415_n310, dp_cluster_3_mult_512_C415_n309,
         dp_cluster_3_mult_512_C415_n308, dp_cluster_3_mult_512_C415_n307,
         dp_cluster_3_mult_512_C415_n306, dp_cluster_3_mult_512_C415_n305,
         dp_cluster_3_mult_512_C415_n304, dp_cluster_3_mult_512_C415_n303,
         dp_cluster_3_mult_512_C415_n302, dp_cluster_3_mult_512_C415_n301,
         dp_cluster_3_mult_512_C415_n300, dp_cluster_3_mult_512_C415_n299,
         dp_cluster_3_mult_512_C415_n298, dp_cluster_3_mult_512_C415_n297,
         dp_cluster_3_mult_512_C415_n296, dp_cluster_3_mult_512_C415_n295,
         dp_cluster_3_mult_512_C415_n294, dp_cluster_3_mult_512_C415_n293,
         dp_cluster_3_mult_512_C415_n292, dp_cluster_3_mult_512_C415_n291,
         dp_cluster_3_mult_512_C415_n290, dp_cluster_3_mult_512_C415_n289,
         dp_cluster_3_mult_512_C415_n288, dp_cluster_3_mult_512_C415_n287,
         dp_cluster_3_mult_512_C415_n286, dp_cluster_3_mult_512_C415_n285,
         dp_cluster_3_mult_512_C415_n284, dp_cluster_3_mult_512_C415_n283,
         dp_cluster_3_mult_512_C415_n282, dp_cluster_3_mult_512_C415_n281,
         dp_cluster_3_mult_512_C415_n280, dp_cluster_3_mult_512_C415_n279,
         dp_cluster_3_mult_512_C415_n278, dp_cluster_3_mult_512_C415_n277,
         dp_cluster_3_mult_512_C415_n275, dp_cluster_3_mult_512_C415_n274,
         dp_cluster_3_mult_512_C415_n273, dp_cluster_3_mult_512_C415_n272,
         dp_cluster_3_mult_512_C415_n271, dp_cluster_3_mult_512_C415_n270,
         dp_cluster_3_mult_512_C415_n269, dp_cluster_3_mult_512_C415_n268,
         dp_cluster_3_mult_512_C415_n267, dp_cluster_3_mult_512_C415_n266,
         dp_cluster_3_mult_512_C415_n264, dp_cluster_3_mult_512_C415_n263,
         dp_cluster_3_mult_512_C415_n262, dp_cluster_3_mult_512_C415_n261,
         dp_cluster_3_mult_512_C415_n260, dp_cluster_3_mult_512_C415_n259,
         dp_cluster_3_mult_512_C415_n258, dp_cluster_3_mult_512_C415_n257,
         dp_cluster_3_mult_512_C415_n256, dp_cluster_3_mult_512_C415_n255,
         dp_cluster_3_mult_512_C415_n254, dp_cluster_3_mult_512_C415_n253,
         dp_cluster_3_mult_512_C415_n252, dp_cluster_3_mult_512_C415_n250,
         dp_cluster_3_mult_512_C415_n249, dp_cluster_3_mult_512_C415_n248,
         dp_cluster_3_mult_512_C415_n247, dp_cluster_3_mult_512_C415_n246,
         dp_cluster_3_mult_512_C415_n245, dp_cluster_3_mult_512_C415_n244,
         dp_cluster_3_mult_512_C415_n243, dp_cluster_3_mult_512_C415_n242,
         dp_cluster_3_mult_512_C415_n241, dp_cluster_3_mult_512_C415_n240,
         dp_cluster_3_mult_512_C415_n239, dp_cluster_3_mult_512_C415_n238,
         dp_cluster_3_mult_512_C415_n237, dp_cluster_3_mult_512_C415_n236,
         dp_cluster_3_mult_512_C415_n235, dp_cluster_3_mult_512_C415_n234,
         dp_cluster_3_mult_512_C415_n233, dp_cluster_3_mult_512_C415_n232,
         dp_cluster_3_mult_512_C415_n231, dp_cluster_3_mult_512_C415_n230,
         dp_cluster_3_mult_512_C415_n229, dp_cluster_3_mult_512_C415_n228,
         dp_cluster_3_mult_512_C415_n227, dp_cluster_3_mult_512_C415_n226,
         dp_cluster_3_mult_512_C415_n225, dp_cluster_3_mult_512_C415_n224,
         dp_cluster_3_mult_512_C415_n223, dp_cluster_3_mult_512_C415_n222,
         dp_cluster_3_mult_512_C415_n221, dp_cluster_3_mult_512_C415_n220,
         dp_cluster_3_mult_512_C415_n219, dp_cluster_3_mult_512_C415_n218,
         dp_cluster_3_mult_512_C415_n217, dp_cluster_3_mult_512_C415_n216,
         dp_cluster_3_mult_512_C415_n215, dp_cluster_3_mult_512_C415_n214,
         dp_cluster_3_mult_512_C415_n213, dp_cluster_3_mult_512_C415_n212,
         dp_cluster_3_mult_512_C415_n211, dp_cluster_3_mult_512_C415_n210,
         dp_cluster_3_mult_512_C415_n209, dp_cluster_3_mult_512_C415_n208,
         dp_cluster_3_mult_512_C415_n207, dp_cluster_3_mult_512_C415_n206,
         dp_cluster_3_mult_512_C415_n205, dp_cluster_3_mult_512_C415_n204,
         dp_cluster_3_mult_512_C415_n203, dp_cluster_3_mult_512_C415_n202,
         dp_cluster_3_mult_512_C415_n201, dp_cluster_3_mult_512_C415_n200,
         dp_cluster_3_mult_512_C415_n199, dp_cluster_3_mult_512_C415_n198,
         dp_cluster_3_mult_512_C415_n197, dp_cluster_3_mult_512_C415_n196,
         dp_cluster_3_mult_512_C415_n195, dp_cluster_3_mult_512_C415_n194,
         dp_cluster_3_mult_512_C415_n193, dp_cluster_3_mult_512_C415_n192,
         dp_cluster_3_mult_512_C415_n191, dp_cluster_3_mult_512_C415_n190,
         dp_cluster_3_mult_512_C415_n189, dp_cluster_3_mult_512_C415_n188,
         dp_cluster_3_mult_512_C415_n187, dp_cluster_3_mult_512_C415_n186,
         dp_cluster_3_mult_512_C415_n185, dp_cluster_3_mult_512_C415_n184,
         dp_cluster_3_mult_512_C415_n183, dp_cluster_3_mult_512_C415_n182,
         dp_cluster_3_mult_512_C415_n181, dp_cluster_3_mult_512_C415_n180,
         dp_cluster_3_mult_512_C415_n179, dp_cluster_3_mult_512_C415_n178,
         dp_cluster_3_mult_512_C415_n177, dp_cluster_3_mult_512_C415_n176,
         dp_cluster_3_mult_512_C415_n175, dp_cluster_3_mult_512_C415_n174,
         dp_cluster_3_mult_512_C415_n173, dp_cluster_3_mult_512_C415_n172,
         dp_cluster_3_mult_512_C415_n171, dp_cluster_3_mult_512_C415_n170,
         dp_cluster_3_mult_512_C415_n169, dp_cluster_3_mult_512_C415_n168,
         dp_cluster_3_mult_512_C415_n167, dp_cluster_3_mult_512_C415_n166,
         dp_cluster_3_mult_512_C415_n165, dp_cluster_3_mult_512_C415_n164,
         dp_cluster_3_mult_512_C415_n163, dp_cluster_3_mult_512_C415_n162,
         dp_cluster_3_mult_512_C415_n161, dp_cluster_3_mult_512_C415_n160,
         dp_cluster_3_mult_512_C415_n159, dp_cluster_3_mult_512_C415_n158,
         dp_cluster_3_mult_512_C415_n157, dp_cluster_3_mult_512_C415_n156,
         dp_cluster_3_mult_512_C415_n155, dp_cluster_3_mult_512_C415_n154,
         dp_cluster_3_mult_512_C415_n153, dp_cluster_3_mult_512_C415_n152,
         dp_cluster_3_mult_512_C415_n150, dp_cluster_3_mult_512_C415_n149,
         dp_cluster_3_mult_512_C415_n148, dp_cluster_3_mult_512_C415_n147,
         dp_cluster_3_mult_512_C415_n146, dp_cluster_3_mult_512_C415_n145,
         dp_cluster_3_mult_512_C415_n144, dp_cluster_3_mult_512_C415_n143,
         dp_cluster_3_mult_512_C415_n142, dp_cluster_3_mult_512_C415_n141,
         dp_cluster_3_mult_512_C415_n140, dp_cluster_3_mult_512_C415_n139,
         dp_cluster_3_mult_512_C415_n138, dp_cluster_3_mult_512_C415_n137,
         dp_cluster_3_mult_512_C415_n136, dp_cluster_3_mult_512_C415_n135,
         dp_cluster_3_mult_512_C415_n134, dp_cluster_3_mult_512_C415_n133,
         dp_cluster_3_mult_512_C415_n132, dp_cluster_3_mult_512_C415_n130,
         dp_cluster_3_mult_512_C415_n129, dp_cluster_3_mult_512_C415_n128,
         dp_cluster_3_mult_512_C415_n127, dp_cluster_3_mult_512_C415_n126,
         dp_cluster_3_mult_512_C415_n125, dp_cluster_3_mult_512_C415_n124,
         dp_cluster_3_mult_512_C415_n123, dp_cluster_3_mult_512_C415_n122,
         dp_cluster_3_mult_512_C415_n121, dp_cluster_3_mult_512_C415_n120,
         dp_cluster_3_mult_512_C415_n119, dp_cluster_3_mult_512_C415_n118,
         dp_cluster_3_mult_512_C415_n117, dp_cluster_3_mult_512_C415_n116,
         dp_cluster_3_mult_512_C415_n115, dp_cluster_3_mult_512_C415_n114,
         dp_cluster_3_mult_512_C415_n112, dp_cluster_3_mult_512_C415_n111,
         dp_cluster_3_mult_512_C415_n110, dp_cluster_3_mult_512_C415_n109,
         dp_cluster_3_mult_512_C415_n108, dp_cluster_3_mult_512_C415_n107,
         dp_cluster_3_mult_512_C415_n106, dp_cluster_3_mult_512_C415_n105,
         dp_cluster_3_mult_512_C415_n104, dp_cluster_3_mult_512_C415_n103,
         dp_cluster_3_mult_512_C415_n102, dp_cluster_3_mult_512_C415_n101,
         dp_cluster_3_mult_512_C415_n100, dp_cluster_3_mult_512_C415_n98,
         dp_cluster_3_mult_512_C415_n97, dp_cluster_3_mult_512_C415_n96,
         dp_cluster_3_mult_512_C415_n95, dp_cluster_3_mult_512_C415_n94,
         dp_cluster_3_mult_512_C415_n93, dp_cluster_3_mult_512_C415_n92,
         dp_cluster_3_mult_512_C415_n91, dp_cluster_3_mult_512_C415_n90,
         dp_cluster_3_mult_512_C415_n89, dp_cluster_3_mult_512_C415_n88,
         dp_cluster_3_mult_512_C415_n86, dp_cluster_3_mult_512_C415_n85,
         dp_cluster_3_mult_512_C415_n84, dp_cluster_3_mult_512_C415_n83,
         dp_cluster_3_mult_512_C415_n82, dp_cluster_3_mult_512_C415_n81,
         dp_cluster_3_mult_512_C415_n80, dp_cluster_3_mult_512_C415_n77,
         dp_cluster_3_mult_512_C415_n76, dp_cluster_3_mult_512_C415_n75,
         dp_cluster_3_mult_512_C415_n74, dp_cluster_3_mult_512_C415_n73,
         dp_cluster_3_mult_512_C415_n72, dp_cluster_3_mult_512_C415_n71,
         dp_cluster_3_mult_512_C415_n70, dp_cluster_3_mult_512_C415_n69,
         dp_cluster_3_mult_512_C415_n68, dp_cluster_3_mult_512_C415_n67,
         dp_cluster_3_mult_512_C415_n66, dp_cluster_3_mult_512_C415_n65,
         dp_cluster_3_mult_512_C415_n64, dp_cluster_3_mult_512_C415_n63,
         dp_cluster_3_mult_512_C415_n62, dp_cluster_3_mult_512_C415_n61,
         dp_cluster_3_mult_512_C415_n60, dp_cluster_3_mult_512_C415_n59,
         dp_cluster_3_mult_512_C415_n58, dp_cluster_3_mult_512_C415_n57,
         dp_cluster_3_mult_512_C415_n56, dp_cluster_3_mult_512_C415_n55,
         dp_cluster_3_mult_512_C415_n54, dp_cluster_3_mult_512_C415_n53,
         dp_cluster_3_mult_512_C415_n52, dp_cluster_3_mult_513_C415_n376,
         dp_cluster_3_mult_513_C415_n375, dp_cluster_3_mult_513_C415_n374,
         dp_cluster_3_mult_513_C415_n373, dp_cluster_3_mult_513_C415_n372,
         dp_cluster_3_mult_513_C415_n371, dp_cluster_3_mult_513_C415_n370,
         dp_cluster_3_mult_513_C415_n369, dp_cluster_3_mult_513_C415_n368,
         dp_cluster_3_mult_513_C415_n367, dp_cluster_3_mult_513_C415_n366,
         dp_cluster_3_mult_513_C415_n365, dp_cluster_3_mult_513_C415_n364,
         dp_cluster_3_mult_513_C415_n363, dp_cluster_3_mult_513_C415_n362,
         dp_cluster_3_mult_513_C415_n361, dp_cluster_3_mult_513_C415_n360,
         dp_cluster_3_mult_513_C415_n359, dp_cluster_3_mult_513_C415_n358,
         dp_cluster_3_mult_513_C415_n357, dp_cluster_3_mult_513_C415_n356,
         dp_cluster_3_mult_513_C415_n355, dp_cluster_3_mult_513_C415_n354,
         dp_cluster_3_mult_513_C415_n353, dp_cluster_3_mult_513_C415_n352,
         dp_cluster_3_mult_513_C415_n351, dp_cluster_3_mult_513_C415_n350,
         dp_cluster_3_mult_513_C415_n349, dp_cluster_3_mult_513_C415_n348,
         dp_cluster_3_mult_513_C415_n347, dp_cluster_3_mult_513_C415_n346,
         dp_cluster_3_mult_513_C415_n345, dp_cluster_3_mult_513_C415_n344,
         dp_cluster_3_mult_513_C415_n343, dp_cluster_3_mult_513_C415_n342,
         dp_cluster_3_mult_513_C415_n341, dp_cluster_3_mult_513_C415_n340,
         dp_cluster_3_mult_513_C415_n339, dp_cluster_3_mult_513_C415_n338,
         dp_cluster_3_mult_513_C415_n337, dp_cluster_3_mult_513_C415_n336,
         dp_cluster_3_mult_513_C415_n335, dp_cluster_3_mult_513_C415_n334,
         dp_cluster_3_mult_513_C415_n333, dp_cluster_3_mult_513_C415_n332,
         dp_cluster_3_mult_513_C415_n331, dp_cluster_3_mult_513_C415_n330,
         dp_cluster_3_mult_513_C415_n329, dp_cluster_3_mult_513_C415_n328,
         dp_cluster_3_mult_513_C415_n327, dp_cluster_3_mult_513_C415_n326,
         dp_cluster_3_mult_513_C415_n325, dp_cluster_3_mult_513_C415_n324,
         dp_cluster_3_mult_513_C415_n323, dp_cluster_3_mult_513_C415_n322,
         dp_cluster_3_mult_513_C415_n321, dp_cluster_3_mult_513_C415_n320,
         dp_cluster_3_mult_513_C415_n319, dp_cluster_3_mult_513_C415_n317,
         dp_cluster_3_mult_513_C415_n316, dp_cluster_3_mult_513_C415_n315,
         dp_cluster_3_mult_513_C415_n314, dp_cluster_3_mult_513_C415_n313,
         dp_cluster_3_mult_513_C415_n312, dp_cluster_3_mult_513_C415_n311,
         dp_cluster_3_mult_513_C415_n310, dp_cluster_3_mult_513_C415_n309,
         dp_cluster_3_mult_513_C415_n308, dp_cluster_3_mult_513_C415_n307,
         dp_cluster_3_mult_513_C415_n306, dp_cluster_3_mult_513_C415_n305,
         dp_cluster_3_mult_513_C415_n304, dp_cluster_3_mult_513_C415_n303,
         dp_cluster_3_mult_513_C415_n302, dp_cluster_3_mult_513_C415_n301,
         dp_cluster_3_mult_513_C415_n300, dp_cluster_3_mult_513_C415_n299,
         dp_cluster_3_mult_513_C415_n298, dp_cluster_3_mult_513_C415_n297,
         dp_cluster_3_mult_513_C415_n296, dp_cluster_3_mult_513_C415_n295,
         dp_cluster_3_mult_513_C415_n294, dp_cluster_3_mult_513_C415_n293,
         dp_cluster_3_mult_513_C415_n292, dp_cluster_3_mult_513_C415_n291,
         dp_cluster_3_mult_513_C415_n290, dp_cluster_3_mult_513_C415_n289,
         dp_cluster_3_mult_513_C415_n288, dp_cluster_3_mult_513_C415_n287,
         dp_cluster_3_mult_513_C415_n286, dp_cluster_3_mult_513_C415_n285,
         dp_cluster_3_mult_513_C415_n284, dp_cluster_3_mult_513_C415_n283,
         dp_cluster_3_mult_513_C415_n282, dp_cluster_3_mult_513_C415_n281,
         dp_cluster_3_mult_513_C415_n280, dp_cluster_3_mult_513_C415_n279,
         dp_cluster_3_mult_513_C415_n278, dp_cluster_3_mult_513_C415_n277,
         dp_cluster_3_mult_513_C415_n275, dp_cluster_3_mult_513_C415_n274,
         dp_cluster_3_mult_513_C415_n273, dp_cluster_3_mult_513_C415_n272,
         dp_cluster_3_mult_513_C415_n271, dp_cluster_3_mult_513_C415_n270,
         dp_cluster_3_mult_513_C415_n269, dp_cluster_3_mult_513_C415_n268,
         dp_cluster_3_mult_513_C415_n267, dp_cluster_3_mult_513_C415_n266,
         dp_cluster_3_mult_513_C415_n264, dp_cluster_3_mult_513_C415_n263,
         dp_cluster_3_mult_513_C415_n262, dp_cluster_3_mult_513_C415_n261,
         dp_cluster_3_mult_513_C415_n260, dp_cluster_3_mult_513_C415_n259,
         dp_cluster_3_mult_513_C415_n258, dp_cluster_3_mult_513_C415_n257,
         dp_cluster_3_mult_513_C415_n256, dp_cluster_3_mult_513_C415_n255,
         dp_cluster_3_mult_513_C415_n254, dp_cluster_3_mult_513_C415_n253,
         dp_cluster_3_mult_513_C415_n252, dp_cluster_3_mult_513_C415_n250,
         dp_cluster_3_mult_513_C415_n249, dp_cluster_3_mult_513_C415_n248,
         dp_cluster_3_mult_513_C415_n247, dp_cluster_3_mult_513_C415_n246,
         dp_cluster_3_mult_513_C415_n245, dp_cluster_3_mult_513_C415_n244,
         dp_cluster_3_mult_513_C415_n243, dp_cluster_3_mult_513_C415_n242,
         dp_cluster_3_mult_513_C415_n241, dp_cluster_3_mult_513_C415_n240,
         dp_cluster_3_mult_513_C415_n239, dp_cluster_3_mult_513_C415_n238,
         dp_cluster_3_mult_513_C415_n237, dp_cluster_3_mult_513_C415_n236,
         dp_cluster_3_mult_513_C415_n235, dp_cluster_3_mult_513_C415_n234,
         dp_cluster_3_mult_513_C415_n233, dp_cluster_3_mult_513_C415_n232,
         dp_cluster_3_mult_513_C415_n231, dp_cluster_3_mult_513_C415_n230,
         dp_cluster_3_mult_513_C415_n229, dp_cluster_3_mult_513_C415_n228,
         dp_cluster_3_mult_513_C415_n227, dp_cluster_3_mult_513_C415_n226,
         dp_cluster_3_mult_513_C415_n225, dp_cluster_3_mult_513_C415_n224,
         dp_cluster_3_mult_513_C415_n223, dp_cluster_3_mult_513_C415_n222,
         dp_cluster_3_mult_513_C415_n221, dp_cluster_3_mult_513_C415_n220,
         dp_cluster_3_mult_513_C415_n219, dp_cluster_3_mult_513_C415_n218,
         dp_cluster_3_mult_513_C415_n217, dp_cluster_3_mult_513_C415_n216,
         dp_cluster_3_mult_513_C415_n215, dp_cluster_3_mult_513_C415_n214,
         dp_cluster_3_mult_513_C415_n213, dp_cluster_3_mult_513_C415_n212,
         dp_cluster_3_mult_513_C415_n211, dp_cluster_3_mult_513_C415_n210,
         dp_cluster_3_mult_513_C415_n209, dp_cluster_3_mult_513_C415_n208,
         dp_cluster_3_mult_513_C415_n207, dp_cluster_3_mult_513_C415_n206,
         dp_cluster_3_mult_513_C415_n205, dp_cluster_3_mult_513_C415_n204,
         dp_cluster_3_mult_513_C415_n203, dp_cluster_3_mult_513_C415_n202,
         dp_cluster_3_mult_513_C415_n201, dp_cluster_3_mult_513_C415_n200,
         dp_cluster_3_mult_513_C415_n199, dp_cluster_3_mult_513_C415_n198,
         dp_cluster_3_mult_513_C415_n197, dp_cluster_3_mult_513_C415_n196,
         dp_cluster_3_mult_513_C415_n195, dp_cluster_3_mult_513_C415_n194,
         dp_cluster_3_mult_513_C415_n193, dp_cluster_3_mult_513_C415_n192,
         dp_cluster_3_mult_513_C415_n191, dp_cluster_3_mult_513_C415_n190,
         dp_cluster_3_mult_513_C415_n189, dp_cluster_3_mult_513_C415_n188,
         dp_cluster_3_mult_513_C415_n187, dp_cluster_3_mult_513_C415_n186,
         dp_cluster_3_mult_513_C415_n185, dp_cluster_3_mult_513_C415_n184,
         dp_cluster_3_mult_513_C415_n183, dp_cluster_3_mult_513_C415_n182,
         dp_cluster_3_mult_513_C415_n181, dp_cluster_3_mult_513_C415_n180,
         dp_cluster_3_mult_513_C415_n179, dp_cluster_3_mult_513_C415_n178,
         dp_cluster_3_mult_513_C415_n177, dp_cluster_3_mult_513_C415_n176,
         dp_cluster_3_mult_513_C415_n175, dp_cluster_3_mult_513_C415_n174,
         dp_cluster_3_mult_513_C415_n173, dp_cluster_3_mult_513_C415_n172,
         dp_cluster_3_mult_513_C415_n171, dp_cluster_3_mult_513_C415_n170,
         dp_cluster_3_mult_513_C415_n169, dp_cluster_3_mult_513_C415_n168,
         dp_cluster_3_mult_513_C415_n167, dp_cluster_3_mult_513_C415_n166,
         dp_cluster_3_mult_513_C415_n165, dp_cluster_3_mult_513_C415_n164,
         dp_cluster_3_mult_513_C415_n163, dp_cluster_3_mult_513_C415_n162,
         dp_cluster_3_mult_513_C415_n161, dp_cluster_3_mult_513_C415_n160,
         dp_cluster_3_mult_513_C415_n159, dp_cluster_3_mult_513_C415_n158,
         dp_cluster_3_mult_513_C415_n157, dp_cluster_3_mult_513_C415_n156,
         dp_cluster_3_mult_513_C415_n155, dp_cluster_3_mult_513_C415_n154,
         dp_cluster_3_mult_513_C415_n153, dp_cluster_3_mult_513_C415_n152,
         dp_cluster_3_mult_513_C415_n150, dp_cluster_3_mult_513_C415_n149,
         dp_cluster_3_mult_513_C415_n148, dp_cluster_3_mult_513_C415_n147,
         dp_cluster_3_mult_513_C415_n146, dp_cluster_3_mult_513_C415_n145,
         dp_cluster_3_mult_513_C415_n144, dp_cluster_3_mult_513_C415_n143,
         dp_cluster_3_mult_513_C415_n142, dp_cluster_3_mult_513_C415_n141,
         dp_cluster_3_mult_513_C415_n140, dp_cluster_3_mult_513_C415_n139,
         dp_cluster_3_mult_513_C415_n138, dp_cluster_3_mult_513_C415_n137,
         dp_cluster_3_mult_513_C415_n136, dp_cluster_3_mult_513_C415_n135,
         dp_cluster_3_mult_513_C415_n134, dp_cluster_3_mult_513_C415_n133,
         dp_cluster_3_mult_513_C415_n132, dp_cluster_3_mult_513_C415_n130,
         dp_cluster_3_mult_513_C415_n129, dp_cluster_3_mult_513_C415_n128,
         dp_cluster_3_mult_513_C415_n127, dp_cluster_3_mult_513_C415_n126,
         dp_cluster_3_mult_513_C415_n125, dp_cluster_3_mult_513_C415_n124,
         dp_cluster_3_mult_513_C415_n123, dp_cluster_3_mult_513_C415_n122,
         dp_cluster_3_mult_513_C415_n121, dp_cluster_3_mult_513_C415_n120,
         dp_cluster_3_mult_513_C415_n119, dp_cluster_3_mult_513_C415_n118,
         dp_cluster_3_mult_513_C415_n117, dp_cluster_3_mult_513_C415_n116,
         dp_cluster_3_mult_513_C415_n115, dp_cluster_3_mult_513_C415_n114,
         dp_cluster_3_mult_513_C415_n112, dp_cluster_3_mult_513_C415_n111,
         dp_cluster_3_mult_513_C415_n110, dp_cluster_3_mult_513_C415_n109,
         dp_cluster_3_mult_513_C415_n108, dp_cluster_3_mult_513_C415_n107,
         dp_cluster_3_mult_513_C415_n106, dp_cluster_3_mult_513_C415_n105,
         dp_cluster_3_mult_513_C415_n104, dp_cluster_3_mult_513_C415_n103,
         dp_cluster_3_mult_513_C415_n102, dp_cluster_3_mult_513_C415_n101,
         dp_cluster_3_mult_513_C415_n100, dp_cluster_3_mult_513_C415_n98,
         dp_cluster_3_mult_513_C415_n97, dp_cluster_3_mult_513_C415_n96,
         dp_cluster_3_mult_513_C415_n95, dp_cluster_3_mult_513_C415_n94,
         dp_cluster_3_mult_513_C415_n93, dp_cluster_3_mult_513_C415_n92,
         dp_cluster_3_mult_513_C415_n91, dp_cluster_3_mult_513_C415_n90,
         dp_cluster_3_mult_513_C415_n89, dp_cluster_3_mult_513_C415_n88,
         dp_cluster_3_mult_513_C415_n86, dp_cluster_3_mult_513_C415_n85,
         dp_cluster_3_mult_513_C415_n84, dp_cluster_3_mult_513_C415_n83,
         dp_cluster_3_mult_513_C415_n82, dp_cluster_3_mult_513_C415_n81,
         dp_cluster_3_mult_513_C415_n80, dp_cluster_3_mult_513_C415_n77,
         dp_cluster_3_mult_513_C415_n76, dp_cluster_3_mult_513_C415_n75,
         dp_cluster_3_mult_513_C415_n74, dp_cluster_3_mult_513_C415_n73,
         dp_cluster_3_mult_513_C415_n72, dp_cluster_3_mult_513_C415_n71,
         dp_cluster_3_mult_513_C415_n70, dp_cluster_3_mult_513_C415_n69,
         dp_cluster_3_mult_513_C415_n68, dp_cluster_3_mult_513_C415_n67,
         dp_cluster_3_mult_513_C415_n66, dp_cluster_3_mult_513_C415_n65,
         dp_cluster_3_mult_513_C415_n64, dp_cluster_3_mult_513_C415_n63,
         dp_cluster_3_mult_513_C415_n62, dp_cluster_3_mult_513_C415_n61,
         dp_cluster_3_mult_513_C415_n60, dp_cluster_3_mult_513_C415_n59,
         dp_cluster_3_mult_513_C415_n58, dp_cluster_3_mult_513_C415_n57,
         dp_cluster_3_mult_513_C415_n56, dp_cluster_3_mult_513_C415_n55,
         dp_cluster_3_mult_513_C415_n54, dp_cluster_3_mult_513_C415_n53,
         dp_cluster_3_mult_513_C415_n52, dp_cluster_2_mult_485_C409_n376,
         dp_cluster_2_mult_485_C409_n375, dp_cluster_2_mult_485_C409_n374,
         dp_cluster_2_mult_485_C409_n373, dp_cluster_2_mult_485_C409_n372,
         dp_cluster_2_mult_485_C409_n371, dp_cluster_2_mult_485_C409_n370,
         dp_cluster_2_mult_485_C409_n369, dp_cluster_2_mult_485_C409_n368,
         dp_cluster_2_mult_485_C409_n367, dp_cluster_2_mult_485_C409_n366,
         dp_cluster_2_mult_485_C409_n365, dp_cluster_2_mult_485_C409_n364,
         dp_cluster_2_mult_485_C409_n363, dp_cluster_2_mult_485_C409_n362,
         dp_cluster_2_mult_485_C409_n361, dp_cluster_2_mult_485_C409_n360,
         dp_cluster_2_mult_485_C409_n359, dp_cluster_2_mult_485_C409_n358,
         dp_cluster_2_mult_485_C409_n357, dp_cluster_2_mult_485_C409_n356,
         dp_cluster_2_mult_485_C409_n355, dp_cluster_2_mult_485_C409_n354,
         dp_cluster_2_mult_485_C409_n353, dp_cluster_2_mult_485_C409_n352,
         dp_cluster_2_mult_485_C409_n351, dp_cluster_2_mult_485_C409_n350,
         dp_cluster_2_mult_485_C409_n349, dp_cluster_2_mult_485_C409_n348,
         dp_cluster_2_mult_485_C409_n347, dp_cluster_2_mult_485_C409_n346,
         dp_cluster_2_mult_485_C409_n345, dp_cluster_2_mult_485_C409_n344,
         dp_cluster_2_mult_485_C409_n343, dp_cluster_2_mult_485_C409_n342,
         dp_cluster_2_mult_485_C409_n341, dp_cluster_2_mult_485_C409_n340,
         dp_cluster_2_mult_485_C409_n339, dp_cluster_2_mult_485_C409_n338,
         dp_cluster_2_mult_485_C409_n337, dp_cluster_2_mult_485_C409_n336,
         dp_cluster_2_mult_485_C409_n335, dp_cluster_2_mult_485_C409_n334,
         dp_cluster_2_mult_485_C409_n333, dp_cluster_2_mult_485_C409_n332,
         dp_cluster_2_mult_485_C409_n331, dp_cluster_2_mult_485_C409_n330,
         dp_cluster_2_mult_485_C409_n329, dp_cluster_2_mult_485_C409_n328,
         dp_cluster_2_mult_485_C409_n327, dp_cluster_2_mult_485_C409_n326,
         dp_cluster_2_mult_485_C409_n325, dp_cluster_2_mult_485_C409_n324,
         dp_cluster_2_mult_485_C409_n323, dp_cluster_2_mult_485_C409_n322,
         dp_cluster_2_mult_485_C409_n321, dp_cluster_2_mult_485_C409_n320,
         dp_cluster_2_mult_485_C409_n319, dp_cluster_2_mult_485_C409_n317,
         dp_cluster_2_mult_485_C409_n316, dp_cluster_2_mult_485_C409_n315,
         dp_cluster_2_mult_485_C409_n314, dp_cluster_2_mult_485_C409_n313,
         dp_cluster_2_mult_485_C409_n312, dp_cluster_2_mult_485_C409_n311,
         dp_cluster_2_mult_485_C409_n310, dp_cluster_2_mult_485_C409_n309,
         dp_cluster_2_mult_485_C409_n308, dp_cluster_2_mult_485_C409_n307,
         dp_cluster_2_mult_485_C409_n306, dp_cluster_2_mult_485_C409_n305,
         dp_cluster_2_mult_485_C409_n304, dp_cluster_2_mult_485_C409_n303,
         dp_cluster_2_mult_485_C409_n302, dp_cluster_2_mult_485_C409_n301,
         dp_cluster_2_mult_485_C409_n300, dp_cluster_2_mult_485_C409_n299,
         dp_cluster_2_mult_485_C409_n298, dp_cluster_2_mult_485_C409_n297,
         dp_cluster_2_mult_485_C409_n296, dp_cluster_2_mult_485_C409_n295,
         dp_cluster_2_mult_485_C409_n294, dp_cluster_2_mult_485_C409_n293,
         dp_cluster_2_mult_485_C409_n292, dp_cluster_2_mult_485_C409_n291,
         dp_cluster_2_mult_485_C409_n290, dp_cluster_2_mult_485_C409_n289,
         dp_cluster_2_mult_485_C409_n288, dp_cluster_2_mult_485_C409_n287,
         dp_cluster_2_mult_485_C409_n286, dp_cluster_2_mult_485_C409_n285,
         dp_cluster_2_mult_485_C409_n284, dp_cluster_2_mult_485_C409_n283,
         dp_cluster_2_mult_485_C409_n282, dp_cluster_2_mult_485_C409_n281,
         dp_cluster_2_mult_485_C409_n280, dp_cluster_2_mult_485_C409_n279,
         dp_cluster_2_mult_485_C409_n278, dp_cluster_2_mult_485_C409_n277,
         dp_cluster_2_mult_485_C409_n275, dp_cluster_2_mult_485_C409_n274,
         dp_cluster_2_mult_485_C409_n273, dp_cluster_2_mult_485_C409_n272,
         dp_cluster_2_mult_485_C409_n271, dp_cluster_2_mult_485_C409_n270,
         dp_cluster_2_mult_485_C409_n269, dp_cluster_2_mult_485_C409_n268,
         dp_cluster_2_mult_485_C409_n267, dp_cluster_2_mult_485_C409_n266,
         dp_cluster_2_mult_485_C409_n264, dp_cluster_2_mult_485_C409_n263,
         dp_cluster_2_mult_485_C409_n262, dp_cluster_2_mult_485_C409_n261,
         dp_cluster_2_mult_485_C409_n260, dp_cluster_2_mult_485_C409_n259,
         dp_cluster_2_mult_485_C409_n258, dp_cluster_2_mult_485_C409_n257,
         dp_cluster_2_mult_485_C409_n256, dp_cluster_2_mult_485_C409_n255,
         dp_cluster_2_mult_485_C409_n254, dp_cluster_2_mult_485_C409_n253,
         dp_cluster_2_mult_485_C409_n252, dp_cluster_2_mult_485_C409_n250,
         dp_cluster_2_mult_485_C409_n249, dp_cluster_2_mult_485_C409_n248,
         dp_cluster_2_mult_485_C409_n247, dp_cluster_2_mult_485_C409_n246,
         dp_cluster_2_mult_485_C409_n245, dp_cluster_2_mult_485_C409_n244,
         dp_cluster_2_mult_485_C409_n243, dp_cluster_2_mult_485_C409_n242,
         dp_cluster_2_mult_485_C409_n241, dp_cluster_2_mult_485_C409_n240,
         dp_cluster_2_mult_485_C409_n239, dp_cluster_2_mult_485_C409_n238,
         dp_cluster_2_mult_485_C409_n237, dp_cluster_2_mult_485_C409_n236,
         dp_cluster_2_mult_485_C409_n235, dp_cluster_2_mult_485_C409_n234,
         dp_cluster_2_mult_485_C409_n233, dp_cluster_2_mult_485_C409_n232,
         dp_cluster_2_mult_485_C409_n231, dp_cluster_2_mult_485_C409_n230,
         dp_cluster_2_mult_485_C409_n229, dp_cluster_2_mult_485_C409_n228,
         dp_cluster_2_mult_485_C409_n227, dp_cluster_2_mult_485_C409_n226,
         dp_cluster_2_mult_485_C409_n225, dp_cluster_2_mult_485_C409_n224,
         dp_cluster_2_mult_485_C409_n223, dp_cluster_2_mult_485_C409_n222,
         dp_cluster_2_mult_485_C409_n221, dp_cluster_2_mult_485_C409_n220,
         dp_cluster_2_mult_485_C409_n219, dp_cluster_2_mult_485_C409_n218,
         dp_cluster_2_mult_485_C409_n217, dp_cluster_2_mult_485_C409_n216,
         dp_cluster_2_mult_485_C409_n215, dp_cluster_2_mult_485_C409_n214,
         dp_cluster_2_mult_485_C409_n213, dp_cluster_2_mult_485_C409_n212,
         dp_cluster_2_mult_485_C409_n211, dp_cluster_2_mult_485_C409_n210,
         dp_cluster_2_mult_485_C409_n209, dp_cluster_2_mult_485_C409_n208,
         dp_cluster_2_mult_485_C409_n207, dp_cluster_2_mult_485_C409_n206,
         dp_cluster_2_mult_485_C409_n205, dp_cluster_2_mult_485_C409_n204,
         dp_cluster_2_mult_485_C409_n203, dp_cluster_2_mult_485_C409_n202,
         dp_cluster_2_mult_485_C409_n201, dp_cluster_2_mult_485_C409_n200,
         dp_cluster_2_mult_485_C409_n199, dp_cluster_2_mult_485_C409_n198,
         dp_cluster_2_mult_485_C409_n197, dp_cluster_2_mult_485_C409_n196,
         dp_cluster_2_mult_485_C409_n195, dp_cluster_2_mult_485_C409_n194,
         dp_cluster_2_mult_485_C409_n193, dp_cluster_2_mult_485_C409_n192,
         dp_cluster_2_mult_485_C409_n191, dp_cluster_2_mult_485_C409_n190,
         dp_cluster_2_mult_485_C409_n189, dp_cluster_2_mult_485_C409_n188,
         dp_cluster_2_mult_485_C409_n187, dp_cluster_2_mult_485_C409_n186,
         dp_cluster_2_mult_485_C409_n185, dp_cluster_2_mult_485_C409_n184,
         dp_cluster_2_mult_485_C409_n183, dp_cluster_2_mult_485_C409_n182,
         dp_cluster_2_mult_485_C409_n181, dp_cluster_2_mult_485_C409_n180,
         dp_cluster_2_mult_485_C409_n179, dp_cluster_2_mult_485_C409_n178,
         dp_cluster_2_mult_485_C409_n177, dp_cluster_2_mult_485_C409_n176,
         dp_cluster_2_mult_485_C409_n175, dp_cluster_2_mult_485_C409_n174,
         dp_cluster_2_mult_485_C409_n173, dp_cluster_2_mult_485_C409_n172,
         dp_cluster_2_mult_485_C409_n171, dp_cluster_2_mult_485_C409_n170,
         dp_cluster_2_mult_485_C409_n169, dp_cluster_2_mult_485_C409_n168,
         dp_cluster_2_mult_485_C409_n167, dp_cluster_2_mult_485_C409_n166,
         dp_cluster_2_mult_485_C409_n165, dp_cluster_2_mult_485_C409_n164,
         dp_cluster_2_mult_485_C409_n163, dp_cluster_2_mult_485_C409_n162,
         dp_cluster_2_mult_485_C409_n161, dp_cluster_2_mult_485_C409_n160,
         dp_cluster_2_mult_485_C409_n159, dp_cluster_2_mult_485_C409_n158,
         dp_cluster_2_mult_485_C409_n157, dp_cluster_2_mult_485_C409_n156,
         dp_cluster_2_mult_485_C409_n155, dp_cluster_2_mult_485_C409_n154,
         dp_cluster_2_mult_485_C409_n153, dp_cluster_2_mult_485_C409_n152,
         dp_cluster_2_mult_485_C409_n150, dp_cluster_2_mult_485_C409_n149,
         dp_cluster_2_mult_485_C409_n148, dp_cluster_2_mult_485_C409_n147,
         dp_cluster_2_mult_485_C409_n146, dp_cluster_2_mult_485_C409_n145,
         dp_cluster_2_mult_485_C409_n144, dp_cluster_2_mult_485_C409_n143,
         dp_cluster_2_mult_485_C409_n142, dp_cluster_2_mult_485_C409_n141,
         dp_cluster_2_mult_485_C409_n140, dp_cluster_2_mult_485_C409_n139,
         dp_cluster_2_mult_485_C409_n138, dp_cluster_2_mult_485_C409_n137,
         dp_cluster_2_mult_485_C409_n136, dp_cluster_2_mult_485_C409_n135,
         dp_cluster_2_mult_485_C409_n134, dp_cluster_2_mult_485_C409_n133,
         dp_cluster_2_mult_485_C409_n132, dp_cluster_2_mult_485_C409_n130,
         dp_cluster_2_mult_485_C409_n129, dp_cluster_2_mult_485_C409_n128,
         dp_cluster_2_mult_485_C409_n127, dp_cluster_2_mult_485_C409_n126,
         dp_cluster_2_mult_485_C409_n125, dp_cluster_2_mult_485_C409_n124,
         dp_cluster_2_mult_485_C409_n123, dp_cluster_2_mult_485_C409_n122,
         dp_cluster_2_mult_485_C409_n121, dp_cluster_2_mult_485_C409_n120,
         dp_cluster_2_mult_485_C409_n119, dp_cluster_2_mult_485_C409_n118,
         dp_cluster_2_mult_485_C409_n117, dp_cluster_2_mult_485_C409_n116,
         dp_cluster_2_mult_485_C409_n115, dp_cluster_2_mult_485_C409_n114,
         dp_cluster_2_mult_485_C409_n112, dp_cluster_2_mult_485_C409_n111,
         dp_cluster_2_mult_485_C409_n110, dp_cluster_2_mult_485_C409_n109,
         dp_cluster_2_mult_485_C409_n108, dp_cluster_2_mult_485_C409_n107,
         dp_cluster_2_mult_485_C409_n106, dp_cluster_2_mult_485_C409_n105,
         dp_cluster_2_mult_485_C409_n104, dp_cluster_2_mult_485_C409_n103,
         dp_cluster_2_mult_485_C409_n102, dp_cluster_2_mult_485_C409_n101,
         dp_cluster_2_mult_485_C409_n100, dp_cluster_2_mult_485_C409_n98,
         dp_cluster_2_mult_485_C409_n97, dp_cluster_2_mult_485_C409_n96,
         dp_cluster_2_mult_485_C409_n95, dp_cluster_2_mult_485_C409_n94,
         dp_cluster_2_mult_485_C409_n93, dp_cluster_2_mult_485_C409_n92,
         dp_cluster_2_mult_485_C409_n91, dp_cluster_2_mult_485_C409_n90,
         dp_cluster_2_mult_485_C409_n89, dp_cluster_2_mult_485_C409_n88,
         dp_cluster_2_mult_485_C409_n86, dp_cluster_2_mult_485_C409_n85,
         dp_cluster_2_mult_485_C409_n84, dp_cluster_2_mult_485_C409_n83,
         dp_cluster_2_mult_485_C409_n82, dp_cluster_2_mult_485_C409_n81,
         dp_cluster_2_mult_485_C409_n80, dp_cluster_2_mult_485_C409_n77,
         dp_cluster_2_mult_485_C409_n76, dp_cluster_2_mult_485_C409_n75,
         dp_cluster_2_mult_485_C409_n74, dp_cluster_2_mult_485_C409_n73,
         dp_cluster_2_mult_485_C409_n72, dp_cluster_2_mult_485_C409_n71,
         dp_cluster_2_mult_485_C409_n70, dp_cluster_2_mult_485_C409_n69,
         dp_cluster_2_mult_485_C409_n68, dp_cluster_2_mult_485_C409_n67,
         dp_cluster_2_mult_485_C409_n66, dp_cluster_2_mult_485_C409_n65,
         dp_cluster_2_mult_485_C409_n64, dp_cluster_2_mult_485_C409_n63,
         dp_cluster_2_mult_485_C409_n62, dp_cluster_2_mult_485_C409_n61,
         dp_cluster_2_mult_485_C409_n60, dp_cluster_2_mult_485_C409_n59,
         dp_cluster_2_mult_485_C409_n58, dp_cluster_2_mult_485_C409_n57,
         dp_cluster_2_mult_485_C409_n56, dp_cluster_2_mult_485_C409_n55,
         dp_cluster_2_mult_485_C409_n54, dp_cluster_2_mult_485_C409_n53,
         dp_cluster_2_mult_485_C409_n52, dp_cluster_2_mult_486_C409_n376,
         dp_cluster_2_mult_486_C409_n375, dp_cluster_2_mult_486_C409_n374,
         dp_cluster_2_mult_486_C409_n373, dp_cluster_2_mult_486_C409_n372,
         dp_cluster_2_mult_486_C409_n371, dp_cluster_2_mult_486_C409_n370,
         dp_cluster_2_mult_486_C409_n369, dp_cluster_2_mult_486_C409_n368,
         dp_cluster_2_mult_486_C409_n367, dp_cluster_2_mult_486_C409_n366,
         dp_cluster_2_mult_486_C409_n365, dp_cluster_2_mult_486_C409_n364,
         dp_cluster_2_mult_486_C409_n363, dp_cluster_2_mult_486_C409_n362,
         dp_cluster_2_mult_486_C409_n361, dp_cluster_2_mult_486_C409_n360,
         dp_cluster_2_mult_486_C409_n359, dp_cluster_2_mult_486_C409_n358,
         dp_cluster_2_mult_486_C409_n357, dp_cluster_2_mult_486_C409_n356,
         dp_cluster_2_mult_486_C409_n355, dp_cluster_2_mult_486_C409_n354,
         dp_cluster_2_mult_486_C409_n353, dp_cluster_2_mult_486_C409_n352,
         dp_cluster_2_mult_486_C409_n351, dp_cluster_2_mult_486_C409_n350,
         dp_cluster_2_mult_486_C409_n349, dp_cluster_2_mult_486_C409_n348,
         dp_cluster_2_mult_486_C409_n347, dp_cluster_2_mult_486_C409_n346,
         dp_cluster_2_mult_486_C409_n345, dp_cluster_2_mult_486_C409_n344,
         dp_cluster_2_mult_486_C409_n343, dp_cluster_2_mult_486_C409_n342,
         dp_cluster_2_mult_486_C409_n341, dp_cluster_2_mult_486_C409_n340,
         dp_cluster_2_mult_486_C409_n339, dp_cluster_2_mult_486_C409_n338,
         dp_cluster_2_mult_486_C409_n337, dp_cluster_2_mult_486_C409_n336,
         dp_cluster_2_mult_486_C409_n335, dp_cluster_2_mult_486_C409_n334,
         dp_cluster_2_mult_486_C409_n333, dp_cluster_2_mult_486_C409_n332,
         dp_cluster_2_mult_486_C409_n331, dp_cluster_2_mult_486_C409_n330,
         dp_cluster_2_mult_486_C409_n329, dp_cluster_2_mult_486_C409_n328,
         dp_cluster_2_mult_486_C409_n327, dp_cluster_2_mult_486_C409_n326,
         dp_cluster_2_mult_486_C409_n325, dp_cluster_2_mult_486_C409_n324,
         dp_cluster_2_mult_486_C409_n323, dp_cluster_2_mult_486_C409_n322,
         dp_cluster_2_mult_486_C409_n321, dp_cluster_2_mult_486_C409_n320,
         dp_cluster_2_mult_486_C409_n319, dp_cluster_2_mult_486_C409_n317,
         dp_cluster_2_mult_486_C409_n316, dp_cluster_2_mult_486_C409_n315,
         dp_cluster_2_mult_486_C409_n314, dp_cluster_2_mult_486_C409_n313,
         dp_cluster_2_mult_486_C409_n312, dp_cluster_2_mult_486_C409_n311,
         dp_cluster_2_mult_486_C409_n310, dp_cluster_2_mult_486_C409_n309,
         dp_cluster_2_mult_486_C409_n308, dp_cluster_2_mult_486_C409_n307,
         dp_cluster_2_mult_486_C409_n306, dp_cluster_2_mult_486_C409_n305,
         dp_cluster_2_mult_486_C409_n304, dp_cluster_2_mult_486_C409_n303,
         dp_cluster_2_mult_486_C409_n302, dp_cluster_2_mult_486_C409_n301,
         dp_cluster_2_mult_486_C409_n300, dp_cluster_2_mult_486_C409_n299,
         dp_cluster_2_mult_486_C409_n298, dp_cluster_2_mult_486_C409_n297,
         dp_cluster_2_mult_486_C409_n296, dp_cluster_2_mult_486_C409_n295,
         dp_cluster_2_mult_486_C409_n294, dp_cluster_2_mult_486_C409_n293,
         dp_cluster_2_mult_486_C409_n292, dp_cluster_2_mult_486_C409_n291,
         dp_cluster_2_mult_486_C409_n290, dp_cluster_2_mult_486_C409_n289,
         dp_cluster_2_mult_486_C409_n288, dp_cluster_2_mult_486_C409_n287,
         dp_cluster_2_mult_486_C409_n286, dp_cluster_2_mult_486_C409_n285,
         dp_cluster_2_mult_486_C409_n284, dp_cluster_2_mult_486_C409_n283,
         dp_cluster_2_mult_486_C409_n282, dp_cluster_2_mult_486_C409_n281,
         dp_cluster_2_mult_486_C409_n280, dp_cluster_2_mult_486_C409_n279,
         dp_cluster_2_mult_486_C409_n278, dp_cluster_2_mult_486_C409_n277,
         dp_cluster_2_mult_486_C409_n275, dp_cluster_2_mult_486_C409_n274,
         dp_cluster_2_mult_486_C409_n273, dp_cluster_2_mult_486_C409_n272,
         dp_cluster_2_mult_486_C409_n271, dp_cluster_2_mult_486_C409_n270,
         dp_cluster_2_mult_486_C409_n269, dp_cluster_2_mult_486_C409_n268,
         dp_cluster_2_mult_486_C409_n267, dp_cluster_2_mult_486_C409_n266,
         dp_cluster_2_mult_486_C409_n264, dp_cluster_2_mult_486_C409_n263,
         dp_cluster_2_mult_486_C409_n262, dp_cluster_2_mult_486_C409_n261,
         dp_cluster_2_mult_486_C409_n260, dp_cluster_2_mult_486_C409_n259,
         dp_cluster_2_mult_486_C409_n258, dp_cluster_2_mult_486_C409_n257,
         dp_cluster_2_mult_486_C409_n256, dp_cluster_2_mult_486_C409_n255,
         dp_cluster_2_mult_486_C409_n254, dp_cluster_2_mult_486_C409_n253,
         dp_cluster_2_mult_486_C409_n252, dp_cluster_2_mult_486_C409_n250,
         dp_cluster_2_mult_486_C409_n249, dp_cluster_2_mult_486_C409_n248,
         dp_cluster_2_mult_486_C409_n247, dp_cluster_2_mult_486_C409_n246,
         dp_cluster_2_mult_486_C409_n245, dp_cluster_2_mult_486_C409_n244,
         dp_cluster_2_mult_486_C409_n243, dp_cluster_2_mult_486_C409_n242,
         dp_cluster_2_mult_486_C409_n241, dp_cluster_2_mult_486_C409_n240,
         dp_cluster_2_mult_486_C409_n239, dp_cluster_2_mult_486_C409_n238,
         dp_cluster_2_mult_486_C409_n237, dp_cluster_2_mult_486_C409_n236,
         dp_cluster_2_mult_486_C409_n235, dp_cluster_2_mult_486_C409_n234,
         dp_cluster_2_mult_486_C409_n233, dp_cluster_2_mult_486_C409_n232,
         dp_cluster_2_mult_486_C409_n231, dp_cluster_2_mult_486_C409_n230,
         dp_cluster_2_mult_486_C409_n229, dp_cluster_2_mult_486_C409_n228,
         dp_cluster_2_mult_486_C409_n227, dp_cluster_2_mult_486_C409_n226,
         dp_cluster_2_mult_486_C409_n225, dp_cluster_2_mult_486_C409_n224,
         dp_cluster_2_mult_486_C409_n223, dp_cluster_2_mult_486_C409_n222,
         dp_cluster_2_mult_486_C409_n221, dp_cluster_2_mult_486_C409_n220,
         dp_cluster_2_mult_486_C409_n219, dp_cluster_2_mult_486_C409_n218,
         dp_cluster_2_mult_486_C409_n217, dp_cluster_2_mult_486_C409_n216,
         dp_cluster_2_mult_486_C409_n215, dp_cluster_2_mult_486_C409_n214,
         dp_cluster_2_mult_486_C409_n213, dp_cluster_2_mult_486_C409_n212,
         dp_cluster_2_mult_486_C409_n211, dp_cluster_2_mult_486_C409_n210,
         dp_cluster_2_mult_486_C409_n209, dp_cluster_2_mult_486_C409_n208,
         dp_cluster_2_mult_486_C409_n207, dp_cluster_2_mult_486_C409_n206,
         dp_cluster_2_mult_486_C409_n205, dp_cluster_2_mult_486_C409_n204,
         dp_cluster_2_mult_486_C409_n203, dp_cluster_2_mult_486_C409_n202,
         dp_cluster_2_mult_486_C409_n201, dp_cluster_2_mult_486_C409_n200,
         dp_cluster_2_mult_486_C409_n199, dp_cluster_2_mult_486_C409_n198,
         dp_cluster_2_mult_486_C409_n197, dp_cluster_2_mult_486_C409_n196,
         dp_cluster_2_mult_486_C409_n195, dp_cluster_2_mult_486_C409_n194,
         dp_cluster_2_mult_486_C409_n193, dp_cluster_2_mult_486_C409_n192,
         dp_cluster_2_mult_486_C409_n191, dp_cluster_2_mult_486_C409_n190,
         dp_cluster_2_mult_486_C409_n189, dp_cluster_2_mult_486_C409_n188,
         dp_cluster_2_mult_486_C409_n187, dp_cluster_2_mult_486_C409_n186,
         dp_cluster_2_mult_486_C409_n185, dp_cluster_2_mult_486_C409_n184,
         dp_cluster_2_mult_486_C409_n183, dp_cluster_2_mult_486_C409_n182,
         dp_cluster_2_mult_486_C409_n181, dp_cluster_2_mult_486_C409_n180,
         dp_cluster_2_mult_486_C409_n179, dp_cluster_2_mult_486_C409_n178,
         dp_cluster_2_mult_486_C409_n177, dp_cluster_2_mult_486_C409_n176,
         dp_cluster_2_mult_486_C409_n175, dp_cluster_2_mult_486_C409_n174,
         dp_cluster_2_mult_486_C409_n173, dp_cluster_2_mult_486_C409_n172,
         dp_cluster_2_mult_486_C409_n171, dp_cluster_2_mult_486_C409_n170,
         dp_cluster_2_mult_486_C409_n169, dp_cluster_2_mult_486_C409_n168,
         dp_cluster_2_mult_486_C409_n167, dp_cluster_2_mult_486_C409_n166,
         dp_cluster_2_mult_486_C409_n165, dp_cluster_2_mult_486_C409_n164,
         dp_cluster_2_mult_486_C409_n163, dp_cluster_2_mult_486_C409_n162,
         dp_cluster_2_mult_486_C409_n161, dp_cluster_2_mult_486_C409_n160,
         dp_cluster_2_mult_486_C409_n159, dp_cluster_2_mult_486_C409_n158,
         dp_cluster_2_mult_486_C409_n157, dp_cluster_2_mult_486_C409_n156,
         dp_cluster_2_mult_486_C409_n155, dp_cluster_2_mult_486_C409_n154,
         dp_cluster_2_mult_486_C409_n153, dp_cluster_2_mult_486_C409_n152,
         dp_cluster_2_mult_486_C409_n150, dp_cluster_2_mult_486_C409_n149,
         dp_cluster_2_mult_486_C409_n148, dp_cluster_2_mult_486_C409_n147,
         dp_cluster_2_mult_486_C409_n146, dp_cluster_2_mult_486_C409_n145,
         dp_cluster_2_mult_486_C409_n144, dp_cluster_2_mult_486_C409_n143,
         dp_cluster_2_mult_486_C409_n142, dp_cluster_2_mult_486_C409_n141,
         dp_cluster_2_mult_486_C409_n140, dp_cluster_2_mult_486_C409_n139,
         dp_cluster_2_mult_486_C409_n138, dp_cluster_2_mult_486_C409_n137,
         dp_cluster_2_mult_486_C409_n136, dp_cluster_2_mult_486_C409_n135,
         dp_cluster_2_mult_486_C409_n134, dp_cluster_2_mult_486_C409_n133,
         dp_cluster_2_mult_486_C409_n132, dp_cluster_2_mult_486_C409_n130,
         dp_cluster_2_mult_486_C409_n129, dp_cluster_2_mult_486_C409_n128,
         dp_cluster_2_mult_486_C409_n127, dp_cluster_2_mult_486_C409_n126,
         dp_cluster_2_mult_486_C409_n125, dp_cluster_2_mult_486_C409_n124,
         dp_cluster_2_mult_486_C409_n123, dp_cluster_2_mult_486_C409_n122,
         dp_cluster_2_mult_486_C409_n121, dp_cluster_2_mult_486_C409_n120,
         dp_cluster_2_mult_486_C409_n119, dp_cluster_2_mult_486_C409_n118,
         dp_cluster_2_mult_486_C409_n117, dp_cluster_2_mult_486_C409_n116,
         dp_cluster_2_mult_486_C409_n115, dp_cluster_2_mult_486_C409_n114,
         dp_cluster_2_mult_486_C409_n112, dp_cluster_2_mult_486_C409_n111,
         dp_cluster_2_mult_486_C409_n110, dp_cluster_2_mult_486_C409_n109,
         dp_cluster_2_mult_486_C409_n108, dp_cluster_2_mult_486_C409_n107,
         dp_cluster_2_mult_486_C409_n106, dp_cluster_2_mult_486_C409_n105,
         dp_cluster_2_mult_486_C409_n104, dp_cluster_2_mult_486_C409_n103,
         dp_cluster_2_mult_486_C409_n102, dp_cluster_2_mult_486_C409_n101,
         dp_cluster_2_mult_486_C409_n100, dp_cluster_2_mult_486_C409_n98,
         dp_cluster_2_mult_486_C409_n97, dp_cluster_2_mult_486_C409_n96,
         dp_cluster_2_mult_486_C409_n95, dp_cluster_2_mult_486_C409_n94,
         dp_cluster_2_mult_486_C409_n93, dp_cluster_2_mult_486_C409_n92,
         dp_cluster_2_mult_486_C409_n91, dp_cluster_2_mult_486_C409_n90,
         dp_cluster_2_mult_486_C409_n89, dp_cluster_2_mult_486_C409_n88,
         dp_cluster_2_mult_486_C409_n86, dp_cluster_2_mult_486_C409_n85,
         dp_cluster_2_mult_486_C409_n84, dp_cluster_2_mult_486_C409_n83,
         dp_cluster_2_mult_486_C409_n82, dp_cluster_2_mult_486_C409_n81,
         dp_cluster_2_mult_486_C409_n80, dp_cluster_2_mult_486_C409_n77,
         dp_cluster_2_mult_486_C409_n76, dp_cluster_2_mult_486_C409_n75,
         dp_cluster_2_mult_486_C409_n74, dp_cluster_2_mult_486_C409_n73,
         dp_cluster_2_mult_486_C409_n72, dp_cluster_2_mult_486_C409_n71,
         dp_cluster_2_mult_486_C409_n70, dp_cluster_2_mult_486_C409_n69,
         dp_cluster_2_mult_486_C409_n68, dp_cluster_2_mult_486_C409_n67,
         dp_cluster_2_mult_486_C409_n66, dp_cluster_2_mult_486_C409_n65,
         dp_cluster_2_mult_486_C409_n64, dp_cluster_2_mult_486_C409_n63,
         dp_cluster_2_mult_486_C409_n62, dp_cluster_2_mult_486_C409_n61,
         dp_cluster_2_mult_486_C409_n60, dp_cluster_2_mult_486_C409_n59,
         dp_cluster_2_mult_486_C409_n58, dp_cluster_2_mult_486_C409_n57,
         dp_cluster_2_mult_486_C409_n56, dp_cluster_2_mult_486_C409_n55,
         dp_cluster_2_mult_486_C409_n54, dp_cluster_2_mult_486_C409_n53,
         dp_cluster_2_mult_486_C409_n52, dp_cluster_1_mult_512_C418_n376,
         dp_cluster_1_mult_512_C418_n375, dp_cluster_1_mult_512_C418_n374,
         dp_cluster_1_mult_512_C418_n373, dp_cluster_1_mult_512_C418_n372,
         dp_cluster_1_mult_512_C418_n371, dp_cluster_1_mult_512_C418_n370,
         dp_cluster_1_mult_512_C418_n369, dp_cluster_1_mult_512_C418_n368,
         dp_cluster_1_mult_512_C418_n367, dp_cluster_1_mult_512_C418_n366,
         dp_cluster_1_mult_512_C418_n365, dp_cluster_1_mult_512_C418_n364,
         dp_cluster_1_mult_512_C418_n363, dp_cluster_1_mult_512_C418_n362,
         dp_cluster_1_mult_512_C418_n361, dp_cluster_1_mult_512_C418_n360,
         dp_cluster_1_mult_512_C418_n359, dp_cluster_1_mult_512_C418_n358,
         dp_cluster_1_mult_512_C418_n357, dp_cluster_1_mult_512_C418_n356,
         dp_cluster_1_mult_512_C418_n355, dp_cluster_1_mult_512_C418_n354,
         dp_cluster_1_mult_512_C418_n353, dp_cluster_1_mult_512_C418_n352,
         dp_cluster_1_mult_512_C418_n351, dp_cluster_1_mult_512_C418_n350,
         dp_cluster_1_mult_512_C418_n349, dp_cluster_1_mult_512_C418_n348,
         dp_cluster_1_mult_512_C418_n347, dp_cluster_1_mult_512_C418_n346,
         dp_cluster_1_mult_512_C418_n345, dp_cluster_1_mult_512_C418_n344,
         dp_cluster_1_mult_512_C418_n343, dp_cluster_1_mult_512_C418_n342,
         dp_cluster_1_mult_512_C418_n341, dp_cluster_1_mult_512_C418_n340,
         dp_cluster_1_mult_512_C418_n339, dp_cluster_1_mult_512_C418_n338,
         dp_cluster_1_mult_512_C418_n337, dp_cluster_1_mult_512_C418_n336,
         dp_cluster_1_mult_512_C418_n335, dp_cluster_1_mult_512_C418_n334,
         dp_cluster_1_mult_512_C418_n333, dp_cluster_1_mult_512_C418_n332,
         dp_cluster_1_mult_512_C418_n331, dp_cluster_1_mult_512_C418_n330,
         dp_cluster_1_mult_512_C418_n329, dp_cluster_1_mult_512_C418_n328,
         dp_cluster_1_mult_512_C418_n327, dp_cluster_1_mult_512_C418_n326,
         dp_cluster_1_mult_512_C418_n325, dp_cluster_1_mult_512_C418_n324,
         dp_cluster_1_mult_512_C418_n323, dp_cluster_1_mult_512_C418_n322,
         dp_cluster_1_mult_512_C418_n321, dp_cluster_1_mult_512_C418_n320,
         dp_cluster_1_mult_512_C418_n319, dp_cluster_1_mult_512_C418_n317,
         dp_cluster_1_mult_512_C418_n316, dp_cluster_1_mult_512_C418_n315,
         dp_cluster_1_mult_512_C418_n314, dp_cluster_1_mult_512_C418_n313,
         dp_cluster_1_mult_512_C418_n312, dp_cluster_1_mult_512_C418_n311,
         dp_cluster_1_mult_512_C418_n310, dp_cluster_1_mult_512_C418_n309,
         dp_cluster_1_mult_512_C418_n308, dp_cluster_1_mult_512_C418_n307,
         dp_cluster_1_mult_512_C418_n306, dp_cluster_1_mult_512_C418_n305,
         dp_cluster_1_mult_512_C418_n304, dp_cluster_1_mult_512_C418_n303,
         dp_cluster_1_mult_512_C418_n302, dp_cluster_1_mult_512_C418_n301,
         dp_cluster_1_mult_512_C418_n300, dp_cluster_1_mult_512_C418_n299,
         dp_cluster_1_mult_512_C418_n298, dp_cluster_1_mult_512_C418_n297,
         dp_cluster_1_mult_512_C418_n296, dp_cluster_1_mult_512_C418_n295,
         dp_cluster_1_mult_512_C418_n294, dp_cluster_1_mult_512_C418_n293,
         dp_cluster_1_mult_512_C418_n292, dp_cluster_1_mult_512_C418_n291,
         dp_cluster_1_mult_512_C418_n290, dp_cluster_1_mult_512_C418_n289,
         dp_cluster_1_mult_512_C418_n288, dp_cluster_1_mult_512_C418_n287,
         dp_cluster_1_mult_512_C418_n286, dp_cluster_1_mult_512_C418_n285,
         dp_cluster_1_mult_512_C418_n284, dp_cluster_1_mult_512_C418_n283,
         dp_cluster_1_mult_512_C418_n282, dp_cluster_1_mult_512_C418_n281,
         dp_cluster_1_mult_512_C418_n280, dp_cluster_1_mult_512_C418_n279,
         dp_cluster_1_mult_512_C418_n278, dp_cluster_1_mult_512_C418_n277,
         dp_cluster_1_mult_512_C418_n275, dp_cluster_1_mult_512_C418_n274,
         dp_cluster_1_mult_512_C418_n273, dp_cluster_1_mult_512_C418_n272,
         dp_cluster_1_mult_512_C418_n271, dp_cluster_1_mult_512_C418_n270,
         dp_cluster_1_mult_512_C418_n269, dp_cluster_1_mult_512_C418_n268,
         dp_cluster_1_mult_512_C418_n267, dp_cluster_1_mult_512_C418_n266,
         dp_cluster_1_mult_512_C418_n264, dp_cluster_1_mult_512_C418_n263,
         dp_cluster_1_mult_512_C418_n262, dp_cluster_1_mult_512_C418_n261,
         dp_cluster_1_mult_512_C418_n260, dp_cluster_1_mult_512_C418_n259,
         dp_cluster_1_mult_512_C418_n258, dp_cluster_1_mult_512_C418_n257,
         dp_cluster_1_mult_512_C418_n256, dp_cluster_1_mult_512_C418_n255,
         dp_cluster_1_mult_512_C418_n254, dp_cluster_1_mult_512_C418_n253,
         dp_cluster_1_mult_512_C418_n252, dp_cluster_1_mult_512_C418_n250,
         dp_cluster_1_mult_512_C418_n249, dp_cluster_1_mult_512_C418_n248,
         dp_cluster_1_mult_512_C418_n247, dp_cluster_1_mult_512_C418_n246,
         dp_cluster_1_mult_512_C418_n245, dp_cluster_1_mult_512_C418_n244,
         dp_cluster_1_mult_512_C418_n243, dp_cluster_1_mult_512_C418_n242,
         dp_cluster_1_mult_512_C418_n241, dp_cluster_1_mult_512_C418_n240,
         dp_cluster_1_mult_512_C418_n239, dp_cluster_1_mult_512_C418_n238,
         dp_cluster_1_mult_512_C418_n237, dp_cluster_1_mult_512_C418_n236,
         dp_cluster_1_mult_512_C418_n235, dp_cluster_1_mult_512_C418_n234,
         dp_cluster_1_mult_512_C418_n233, dp_cluster_1_mult_512_C418_n232,
         dp_cluster_1_mult_512_C418_n231, dp_cluster_1_mult_512_C418_n230,
         dp_cluster_1_mult_512_C418_n229, dp_cluster_1_mult_512_C418_n228,
         dp_cluster_1_mult_512_C418_n227, dp_cluster_1_mult_512_C418_n226,
         dp_cluster_1_mult_512_C418_n225, dp_cluster_1_mult_512_C418_n224,
         dp_cluster_1_mult_512_C418_n223, dp_cluster_1_mult_512_C418_n222,
         dp_cluster_1_mult_512_C418_n221, dp_cluster_1_mult_512_C418_n220,
         dp_cluster_1_mult_512_C418_n219, dp_cluster_1_mult_512_C418_n218,
         dp_cluster_1_mult_512_C418_n217, dp_cluster_1_mult_512_C418_n216,
         dp_cluster_1_mult_512_C418_n215, dp_cluster_1_mult_512_C418_n214,
         dp_cluster_1_mult_512_C418_n213, dp_cluster_1_mult_512_C418_n212,
         dp_cluster_1_mult_512_C418_n211, dp_cluster_1_mult_512_C418_n210,
         dp_cluster_1_mult_512_C418_n209, dp_cluster_1_mult_512_C418_n208,
         dp_cluster_1_mult_512_C418_n207, dp_cluster_1_mult_512_C418_n206,
         dp_cluster_1_mult_512_C418_n205, dp_cluster_1_mult_512_C418_n204,
         dp_cluster_1_mult_512_C418_n203, dp_cluster_1_mult_512_C418_n202,
         dp_cluster_1_mult_512_C418_n201, dp_cluster_1_mult_512_C418_n200,
         dp_cluster_1_mult_512_C418_n199, dp_cluster_1_mult_512_C418_n198,
         dp_cluster_1_mult_512_C418_n197, dp_cluster_1_mult_512_C418_n196,
         dp_cluster_1_mult_512_C418_n195, dp_cluster_1_mult_512_C418_n194,
         dp_cluster_1_mult_512_C418_n193, dp_cluster_1_mult_512_C418_n192,
         dp_cluster_1_mult_512_C418_n191, dp_cluster_1_mult_512_C418_n190,
         dp_cluster_1_mult_512_C418_n189, dp_cluster_1_mult_512_C418_n188,
         dp_cluster_1_mult_512_C418_n187, dp_cluster_1_mult_512_C418_n186,
         dp_cluster_1_mult_512_C418_n185, dp_cluster_1_mult_512_C418_n184,
         dp_cluster_1_mult_512_C418_n183, dp_cluster_1_mult_512_C418_n182,
         dp_cluster_1_mult_512_C418_n181, dp_cluster_1_mult_512_C418_n180,
         dp_cluster_1_mult_512_C418_n179, dp_cluster_1_mult_512_C418_n178,
         dp_cluster_1_mult_512_C418_n177, dp_cluster_1_mult_512_C418_n176,
         dp_cluster_1_mult_512_C418_n175, dp_cluster_1_mult_512_C418_n174,
         dp_cluster_1_mult_512_C418_n173, dp_cluster_1_mult_512_C418_n172,
         dp_cluster_1_mult_512_C418_n171, dp_cluster_1_mult_512_C418_n170,
         dp_cluster_1_mult_512_C418_n169, dp_cluster_1_mult_512_C418_n168,
         dp_cluster_1_mult_512_C418_n167, dp_cluster_1_mult_512_C418_n166,
         dp_cluster_1_mult_512_C418_n165, dp_cluster_1_mult_512_C418_n164,
         dp_cluster_1_mult_512_C418_n163, dp_cluster_1_mult_512_C418_n162,
         dp_cluster_1_mult_512_C418_n161, dp_cluster_1_mult_512_C418_n160,
         dp_cluster_1_mult_512_C418_n159, dp_cluster_1_mult_512_C418_n158,
         dp_cluster_1_mult_512_C418_n157, dp_cluster_1_mult_512_C418_n156,
         dp_cluster_1_mult_512_C418_n155, dp_cluster_1_mult_512_C418_n154,
         dp_cluster_1_mult_512_C418_n153, dp_cluster_1_mult_512_C418_n152,
         dp_cluster_1_mult_512_C418_n150, dp_cluster_1_mult_512_C418_n149,
         dp_cluster_1_mult_512_C418_n148, dp_cluster_1_mult_512_C418_n147,
         dp_cluster_1_mult_512_C418_n146, dp_cluster_1_mult_512_C418_n145,
         dp_cluster_1_mult_512_C418_n144, dp_cluster_1_mult_512_C418_n143,
         dp_cluster_1_mult_512_C418_n142, dp_cluster_1_mult_512_C418_n141,
         dp_cluster_1_mult_512_C418_n140, dp_cluster_1_mult_512_C418_n139,
         dp_cluster_1_mult_512_C418_n138, dp_cluster_1_mult_512_C418_n137,
         dp_cluster_1_mult_512_C418_n136, dp_cluster_1_mult_512_C418_n135,
         dp_cluster_1_mult_512_C418_n134, dp_cluster_1_mult_512_C418_n133,
         dp_cluster_1_mult_512_C418_n132, dp_cluster_1_mult_512_C418_n130,
         dp_cluster_1_mult_512_C418_n129, dp_cluster_1_mult_512_C418_n128,
         dp_cluster_1_mult_512_C418_n127, dp_cluster_1_mult_512_C418_n126,
         dp_cluster_1_mult_512_C418_n125, dp_cluster_1_mult_512_C418_n124,
         dp_cluster_1_mult_512_C418_n123, dp_cluster_1_mult_512_C418_n122,
         dp_cluster_1_mult_512_C418_n121, dp_cluster_1_mult_512_C418_n120,
         dp_cluster_1_mult_512_C418_n119, dp_cluster_1_mult_512_C418_n118,
         dp_cluster_1_mult_512_C418_n117, dp_cluster_1_mult_512_C418_n116,
         dp_cluster_1_mult_512_C418_n115, dp_cluster_1_mult_512_C418_n114,
         dp_cluster_1_mult_512_C418_n112, dp_cluster_1_mult_512_C418_n111,
         dp_cluster_1_mult_512_C418_n110, dp_cluster_1_mult_512_C418_n109,
         dp_cluster_1_mult_512_C418_n108, dp_cluster_1_mult_512_C418_n107,
         dp_cluster_1_mult_512_C418_n106, dp_cluster_1_mult_512_C418_n105,
         dp_cluster_1_mult_512_C418_n104, dp_cluster_1_mult_512_C418_n103,
         dp_cluster_1_mult_512_C418_n102, dp_cluster_1_mult_512_C418_n101,
         dp_cluster_1_mult_512_C418_n100, dp_cluster_1_mult_512_C418_n98,
         dp_cluster_1_mult_512_C418_n97, dp_cluster_1_mult_512_C418_n96,
         dp_cluster_1_mult_512_C418_n95, dp_cluster_1_mult_512_C418_n94,
         dp_cluster_1_mult_512_C418_n93, dp_cluster_1_mult_512_C418_n92,
         dp_cluster_1_mult_512_C418_n91, dp_cluster_1_mult_512_C418_n90,
         dp_cluster_1_mult_512_C418_n89, dp_cluster_1_mult_512_C418_n88,
         dp_cluster_1_mult_512_C418_n86, dp_cluster_1_mult_512_C418_n85,
         dp_cluster_1_mult_512_C418_n84, dp_cluster_1_mult_512_C418_n83,
         dp_cluster_1_mult_512_C418_n82, dp_cluster_1_mult_512_C418_n81,
         dp_cluster_1_mult_512_C418_n80, dp_cluster_1_mult_512_C418_n77,
         dp_cluster_1_mult_512_C418_n76, dp_cluster_1_mult_512_C418_n75,
         dp_cluster_1_mult_512_C418_n74, dp_cluster_1_mult_512_C418_n73,
         dp_cluster_1_mult_512_C418_n72, dp_cluster_1_mult_512_C418_n71,
         dp_cluster_1_mult_512_C418_n70, dp_cluster_1_mult_512_C418_n69,
         dp_cluster_1_mult_512_C418_n68, dp_cluster_1_mult_512_C418_n67,
         dp_cluster_1_mult_512_C418_n66, dp_cluster_1_mult_512_C418_n65,
         dp_cluster_1_mult_512_C418_n64, dp_cluster_1_mult_512_C418_n63,
         dp_cluster_1_mult_512_C418_n62, dp_cluster_1_mult_512_C418_n61,
         dp_cluster_1_mult_512_C418_n60, dp_cluster_1_mult_512_C418_n59,
         dp_cluster_1_mult_512_C418_n58, dp_cluster_1_mult_512_C418_n57,
         dp_cluster_1_mult_512_C418_n56, dp_cluster_1_mult_512_C418_n55,
         dp_cluster_1_mult_512_C418_n54, dp_cluster_1_mult_512_C418_n53,
         dp_cluster_1_mult_512_C418_n52, dp_cluster_1_mult_513_C418_n376,
         dp_cluster_1_mult_513_C418_n375, dp_cluster_1_mult_513_C418_n374,
         dp_cluster_1_mult_513_C418_n373, dp_cluster_1_mult_513_C418_n372,
         dp_cluster_1_mult_513_C418_n371, dp_cluster_1_mult_513_C418_n370,
         dp_cluster_1_mult_513_C418_n369, dp_cluster_1_mult_513_C418_n368,
         dp_cluster_1_mult_513_C418_n367, dp_cluster_1_mult_513_C418_n366,
         dp_cluster_1_mult_513_C418_n365, dp_cluster_1_mult_513_C418_n364,
         dp_cluster_1_mult_513_C418_n363, dp_cluster_1_mult_513_C418_n362,
         dp_cluster_1_mult_513_C418_n361, dp_cluster_1_mult_513_C418_n360,
         dp_cluster_1_mult_513_C418_n359, dp_cluster_1_mult_513_C418_n358,
         dp_cluster_1_mult_513_C418_n357, dp_cluster_1_mult_513_C418_n356,
         dp_cluster_1_mult_513_C418_n355, dp_cluster_1_mult_513_C418_n354,
         dp_cluster_1_mult_513_C418_n353, dp_cluster_1_mult_513_C418_n352,
         dp_cluster_1_mult_513_C418_n351, dp_cluster_1_mult_513_C418_n350,
         dp_cluster_1_mult_513_C418_n349, dp_cluster_1_mult_513_C418_n348,
         dp_cluster_1_mult_513_C418_n347, dp_cluster_1_mult_513_C418_n346,
         dp_cluster_1_mult_513_C418_n345, dp_cluster_1_mult_513_C418_n344,
         dp_cluster_1_mult_513_C418_n343, dp_cluster_1_mult_513_C418_n342,
         dp_cluster_1_mult_513_C418_n341, dp_cluster_1_mult_513_C418_n340,
         dp_cluster_1_mult_513_C418_n339, dp_cluster_1_mult_513_C418_n338,
         dp_cluster_1_mult_513_C418_n337, dp_cluster_1_mult_513_C418_n336,
         dp_cluster_1_mult_513_C418_n335, dp_cluster_1_mult_513_C418_n334,
         dp_cluster_1_mult_513_C418_n333, dp_cluster_1_mult_513_C418_n332,
         dp_cluster_1_mult_513_C418_n331, dp_cluster_1_mult_513_C418_n330,
         dp_cluster_1_mult_513_C418_n329, dp_cluster_1_mult_513_C418_n328,
         dp_cluster_1_mult_513_C418_n327, dp_cluster_1_mult_513_C418_n326,
         dp_cluster_1_mult_513_C418_n325, dp_cluster_1_mult_513_C418_n324,
         dp_cluster_1_mult_513_C418_n323, dp_cluster_1_mult_513_C418_n322,
         dp_cluster_1_mult_513_C418_n321, dp_cluster_1_mult_513_C418_n320,
         dp_cluster_1_mult_513_C418_n319, dp_cluster_1_mult_513_C418_n317,
         dp_cluster_1_mult_513_C418_n316, dp_cluster_1_mult_513_C418_n315,
         dp_cluster_1_mult_513_C418_n314, dp_cluster_1_mult_513_C418_n313,
         dp_cluster_1_mult_513_C418_n312, dp_cluster_1_mult_513_C418_n311,
         dp_cluster_1_mult_513_C418_n310, dp_cluster_1_mult_513_C418_n309,
         dp_cluster_1_mult_513_C418_n308, dp_cluster_1_mult_513_C418_n307,
         dp_cluster_1_mult_513_C418_n306, dp_cluster_1_mult_513_C418_n305,
         dp_cluster_1_mult_513_C418_n304, dp_cluster_1_mult_513_C418_n303,
         dp_cluster_1_mult_513_C418_n302, dp_cluster_1_mult_513_C418_n301,
         dp_cluster_1_mult_513_C418_n300, dp_cluster_1_mult_513_C418_n299,
         dp_cluster_1_mult_513_C418_n298, dp_cluster_1_mult_513_C418_n297,
         dp_cluster_1_mult_513_C418_n296, dp_cluster_1_mult_513_C418_n295,
         dp_cluster_1_mult_513_C418_n294, dp_cluster_1_mult_513_C418_n293,
         dp_cluster_1_mult_513_C418_n292, dp_cluster_1_mult_513_C418_n291,
         dp_cluster_1_mult_513_C418_n290, dp_cluster_1_mult_513_C418_n289,
         dp_cluster_1_mult_513_C418_n288, dp_cluster_1_mult_513_C418_n287,
         dp_cluster_1_mult_513_C418_n286, dp_cluster_1_mult_513_C418_n285,
         dp_cluster_1_mult_513_C418_n284, dp_cluster_1_mult_513_C418_n283,
         dp_cluster_1_mult_513_C418_n282, dp_cluster_1_mult_513_C418_n281,
         dp_cluster_1_mult_513_C418_n280, dp_cluster_1_mult_513_C418_n279,
         dp_cluster_1_mult_513_C418_n278, dp_cluster_1_mult_513_C418_n277,
         dp_cluster_1_mult_513_C418_n275, dp_cluster_1_mult_513_C418_n274,
         dp_cluster_1_mult_513_C418_n273, dp_cluster_1_mult_513_C418_n272,
         dp_cluster_1_mult_513_C418_n271, dp_cluster_1_mult_513_C418_n270,
         dp_cluster_1_mult_513_C418_n269, dp_cluster_1_mult_513_C418_n268,
         dp_cluster_1_mult_513_C418_n267, dp_cluster_1_mult_513_C418_n266,
         dp_cluster_1_mult_513_C418_n264, dp_cluster_1_mult_513_C418_n263,
         dp_cluster_1_mult_513_C418_n262, dp_cluster_1_mult_513_C418_n261,
         dp_cluster_1_mult_513_C418_n260, dp_cluster_1_mult_513_C418_n259,
         dp_cluster_1_mult_513_C418_n258, dp_cluster_1_mult_513_C418_n257,
         dp_cluster_1_mult_513_C418_n256, dp_cluster_1_mult_513_C418_n255,
         dp_cluster_1_mult_513_C418_n254, dp_cluster_1_mult_513_C418_n253,
         dp_cluster_1_mult_513_C418_n252, dp_cluster_1_mult_513_C418_n250,
         dp_cluster_1_mult_513_C418_n249, dp_cluster_1_mult_513_C418_n248,
         dp_cluster_1_mult_513_C418_n247, dp_cluster_1_mult_513_C418_n246,
         dp_cluster_1_mult_513_C418_n245, dp_cluster_1_mult_513_C418_n244,
         dp_cluster_1_mult_513_C418_n243, dp_cluster_1_mult_513_C418_n242,
         dp_cluster_1_mult_513_C418_n241, dp_cluster_1_mult_513_C418_n240,
         dp_cluster_1_mult_513_C418_n239, dp_cluster_1_mult_513_C418_n238,
         dp_cluster_1_mult_513_C418_n237, dp_cluster_1_mult_513_C418_n236,
         dp_cluster_1_mult_513_C418_n235, dp_cluster_1_mult_513_C418_n234,
         dp_cluster_1_mult_513_C418_n233, dp_cluster_1_mult_513_C418_n232,
         dp_cluster_1_mult_513_C418_n231, dp_cluster_1_mult_513_C418_n230,
         dp_cluster_1_mult_513_C418_n229, dp_cluster_1_mult_513_C418_n228,
         dp_cluster_1_mult_513_C418_n227, dp_cluster_1_mult_513_C418_n226,
         dp_cluster_1_mult_513_C418_n225, dp_cluster_1_mult_513_C418_n224,
         dp_cluster_1_mult_513_C418_n223, dp_cluster_1_mult_513_C418_n222,
         dp_cluster_1_mult_513_C418_n221, dp_cluster_1_mult_513_C418_n220,
         dp_cluster_1_mult_513_C418_n219, dp_cluster_1_mult_513_C418_n218,
         dp_cluster_1_mult_513_C418_n217, dp_cluster_1_mult_513_C418_n216,
         dp_cluster_1_mult_513_C418_n215, dp_cluster_1_mult_513_C418_n214,
         dp_cluster_1_mult_513_C418_n213, dp_cluster_1_mult_513_C418_n212,
         dp_cluster_1_mult_513_C418_n211, dp_cluster_1_mult_513_C418_n210,
         dp_cluster_1_mult_513_C418_n209, dp_cluster_1_mult_513_C418_n208,
         dp_cluster_1_mult_513_C418_n207, dp_cluster_1_mult_513_C418_n206,
         dp_cluster_1_mult_513_C418_n205, dp_cluster_1_mult_513_C418_n204,
         dp_cluster_1_mult_513_C418_n203, dp_cluster_1_mult_513_C418_n202,
         dp_cluster_1_mult_513_C418_n201, dp_cluster_1_mult_513_C418_n200,
         dp_cluster_1_mult_513_C418_n199, dp_cluster_1_mult_513_C418_n198,
         dp_cluster_1_mult_513_C418_n197, dp_cluster_1_mult_513_C418_n196,
         dp_cluster_1_mult_513_C418_n195, dp_cluster_1_mult_513_C418_n194,
         dp_cluster_1_mult_513_C418_n193, dp_cluster_1_mult_513_C418_n192,
         dp_cluster_1_mult_513_C418_n191, dp_cluster_1_mult_513_C418_n190,
         dp_cluster_1_mult_513_C418_n189, dp_cluster_1_mult_513_C418_n188,
         dp_cluster_1_mult_513_C418_n187, dp_cluster_1_mult_513_C418_n186,
         dp_cluster_1_mult_513_C418_n185, dp_cluster_1_mult_513_C418_n184,
         dp_cluster_1_mult_513_C418_n183, dp_cluster_1_mult_513_C418_n182,
         dp_cluster_1_mult_513_C418_n181, dp_cluster_1_mult_513_C418_n180,
         dp_cluster_1_mult_513_C418_n179, dp_cluster_1_mult_513_C418_n178,
         dp_cluster_1_mult_513_C418_n177, dp_cluster_1_mult_513_C418_n176,
         dp_cluster_1_mult_513_C418_n175, dp_cluster_1_mult_513_C418_n174,
         dp_cluster_1_mult_513_C418_n173, dp_cluster_1_mult_513_C418_n172,
         dp_cluster_1_mult_513_C418_n171, dp_cluster_1_mult_513_C418_n170,
         dp_cluster_1_mult_513_C418_n169, dp_cluster_1_mult_513_C418_n168,
         dp_cluster_1_mult_513_C418_n167, dp_cluster_1_mult_513_C418_n166,
         dp_cluster_1_mult_513_C418_n165, dp_cluster_1_mult_513_C418_n164,
         dp_cluster_1_mult_513_C418_n163, dp_cluster_1_mult_513_C418_n162,
         dp_cluster_1_mult_513_C418_n161, dp_cluster_1_mult_513_C418_n160,
         dp_cluster_1_mult_513_C418_n159, dp_cluster_1_mult_513_C418_n158,
         dp_cluster_1_mult_513_C418_n157, dp_cluster_1_mult_513_C418_n156,
         dp_cluster_1_mult_513_C418_n155, dp_cluster_1_mult_513_C418_n154,
         dp_cluster_1_mult_513_C418_n153, dp_cluster_1_mult_513_C418_n152,
         dp_cluster_1_mult_513_C418_n150, dp_cluster_1_mult_513_C418_n149,
         dp_cluster_1_mult_513_C418_n148, dp_cluster_1_mult_513_C418_n147,
         dp_cluster_1_mult_513_C418_n146, dp_cluster_1_mult_513_C418_n145,
         dp_cluster_1_mult_513_C418_n144, dp_cluster_1_mult_513_C418_n143,
         dp_cluster_1_mult_513_C418_n142, dp_cluster_1_mult_513_C418_n141,
         dp_cluster_1_mult_513_C418_n140, dp_cluster_1_mult_513_C418_n139,
         dp_cluster_1_mult_513_C418_n138, dp_cluster_1_mult_513_C418_n137,
         dp_cluster_1_mult_513_C418_n136, dp_cluster_1_mult_513_C418_n135,
         dp_cluster_1_mult_513_C418_n134, dp_cluster_1_mult_513_C418_n133,
         dp_cluster_1_mult_513_C418_n132, dp_cluster_1_mult_513_C418_n130,
         dp_cluster_1_mult_513_C418_n129, dp_cluster_1_mult_513_C418_n128,
         dp_cluster_1_mult_513_C418_n127, dp_cluster_1_mult_513_C418_n126,
         dp_cluster_1_mult_513_C418_n125, dp_cluster_1_mult_513_C418_n124,
         dp_cluster_1_mult_513_C418_n123, dp_cluster_1_mult_513_C418_n122,
         dp_cluster_1_mult_513_C418_n121, dp_cluster_1_mult_513_C418_n120,
         dp_cluster_1_mult_513_C418_n119, dp_cluster_1_mult_513_C418_n118,
         dp_cluster_1_mult_513_C418_n117, dp_cluster_1_mult_513_C418_n116,
         dp_cluster_1_mult_513_C418_n115, dp_cluster_1_mult_513_C418_n114,
         dp_cluster_1_mult_513_C418_n112, dp_cluster_1_mult_513_C418_n111,
         dp_cluster_1_mult_513_C418_n110, dp_cluster_1_mult_513_C418_n109,
         dp_cluster_1_mult_513_C418_n108, dp_cluster_1_mult_513_C418_n107,
         dp_cluster_1_mult_513_C418_n106, dp_cluster_1_mult_513_C418_n105,
         dp_cluster_1_mult_513_C418_n104, dp_cluster_1_mult_513_C418_n103,
         dp_cluster_1_mult_513_C418_n102, dp_cluster_1_mult_513_C418_n101,
         dp_cluster_1_mult_513_C418_n100, dp_cluster_1_mult_513_C418_n98,
         dp_cluster_1_mult_513_C418_n97, dp_cluster_1_mult_513_C418_n96,
         dp_cluster_1_mult_513_C418_n95, dp_cluster_1_mult_513_C418_n94,
         dp_cluster_1_mult_513_C418_n93, dp_cluster_1_mult_513_C418_n92,
         dp_cluster_1_mult_513_C418_n91, dp_cluster_1_mult_513_C418_n90,
         dp_cluster_1_mult_513_C418_n89, dp_cluster_1_mult_513_C418_n88,
         dp_cluster_1_mult_513_C418_n86, dp_cluster_1_mult_513_C418_n85,
         dp_cluster_1_mult_513_C418_n84, dp_cluster_1_mult_513_C418_n83,
         dp_cluster_1_mult_513_C418_n82, dp_cluster_1_mult_513_C418_n81,
         dp_cluster_1_mult_513_C418_n80, dp_cluster_1_mult_513_C418_n77,
         dp_cluster_1_mult_513_C418_n76, dp_cluster_1_mult_513_C418_n75,
         dp_cluster_1_mult_513_C418_n74, dp_cluster_1_mult_513_C418_n73,
         dp_cluster_1_mult_513_C418_n72, dp_cluster_1_mult_513_C418_n71,
         dp_cluster_1_mult_513_C418_n70, dp_cluster_1_mult_513_C418_n69,
         dp_cluster_1_mult_513_C418_n68, dp_cluster_1_mult_513_C418_n67,
         dp_cluster_1_mult_513_C418_n66, dp_cluster_1_mult_513_C418_n65,
         dp_cluster_1_mult_513_C418_n64, dp_cluster_1_mult_513_C418_n63,
         dp_cluster_1_mult_513_C418_n62, dp_cluster_1_mult_513_C418_n61,
         dp_cluster_1_mult_513_C418_n60, dp_cluster_1_mult_513_C418_n59,
         dp_cluster_1_mult_513_C418_n58, dp_cluster_1_mult_513_C418_n57,
         dp_cluster_1_mult_513_C418_n56, dp_cluster_1_mult_513_C418_n55,
         dp_cluster_1_mult_513_C418_n54, dp_cluster_1_mult_513_C418_n53,
         dp_cluster_1_mult_513_C418_n52, dp_cluster_0_mult_485_C412_n376,
         dp_cluster_0_mult_485_C412_n375, dp_cluster_0_mult_485_C412_n374,
         dp_cluster_0_mult_485_C412_n373, dp_cluster_0_mult_485_C412_n372,
         dp_cluster_0_mult_485_C412_n371, dp_cluster_0_mult_485_C412_n370,
         dp_cluster_0_mult_485_C412_n369, dp_cluster_0_mult_485_C412_n368,
         dp_cluster_0_mult_485_C412_n367, dp_cluster_0_mult_485_C412_n366,
         dp_cluster_0_mult_485_C412_n365, dp_cluster_0_mult_485_C412_n364,
         dp_cluster_0_mult_485_C412_n363, dp_cluster_0_mult_485_C412_n362,
         dp_cluster_0_mult_485_C412_n361, dp_cluster_0_mult_485_C412_n360,
         dp_cluster_0_mult_485_C412_n359, dp_cluster_0_mult_485_C412_n358,
         dp_cluster_0_mult_485_C412_n357, dp_cluster_0_mult_485_C412_n356,
         dp_cluster_0_mult_485_C412_n355, dp_cluster_0_mult_485_C412_n354,
         dp_cluster_0_mult_485_C412_n353, dp_cluster_0_mult_485_C412_n352,
         dp_cluster_0_mult_485_C412_n351, dp_cluster_0_mult_485_C412_n350,
         dp_cluster_0_mult_485_C412_n349, dp_cluster_0_mult_485_C412_n348,
         dp_cluster_0_mult_485_C412_n347, dp_cluster_0_mult_485_C412_n346,
         dp_cluster_0_mult_485_C412_n345, dp_cluster_0_mult_485_C412_n344,
         dp_cluster_0_mult_485_C412_n343, dp_cluster_0_mult_485_C412_n342,
         dp_cluster_0_mult_485_C412_n341, dp_cluster_0_mult_485_C412_n340,
         dp_cluster_0_mult_485_C412_n339, dp_cluster_0_mult_485_C412_n338,
         dp_cluster_0_mult_485_C412_n337, dp_cluster_0_mult_485_C412_n336,
         dp_cluster_0_mult_485_C412_n335, dp_cluster_0_mult_485_C412_n334,
         dp_cluster_0_mult_485_C412_n333, dp_cluster_0_mult_485_C412_n332,
         dp_cluster_0_mult_485_C412_n331, dp_cluster_0_mult_485_C412_n330,
         dp_cluster_0_mult_485_C412_n329, dp_cluster_0_mult_485_C412_n328,
         dp_cluster_0_mult_485_C412_n327, dp_cluster_0_mult_485_C412_n326,
         dp_cluster_0_mult_485_C412_n325, dp_cluster_0_mult_485_C412_n324,
         dp_cluster_0_mult_485_C412_n323, dp_cluster_0_mult_485_C412_n322,
         dp_cluster_0_mult_485_C412_n321, dp_cluster_0_mult_485_C412_n320,
         dp_cluster_0_mult_485_C412_n319, dp_cluster_0_mult_485_C412_n317,
         dp_cluster_0_mult_485_C412_n316, dp_cluster_0_mult_485_C412_n315,
         dp_cluster_0_mult_485_C412_n314, dp_cluster_0_mult_485_C412_n313,
         dp_cluster_0_mult_485_C412_n312, dp_cluster_0_mult_485_C412_n311,
         dp_cluster_0_mult_485_C412_n310, dp_cluster_0_mult_485_C412_n309,
         dp_cluster_0_mult_485_C412_n308, dp_cluster_0_mult_485_C412_n307,
         dp_cluster_0_mult_485_C412_n306, dp_cluster_0_mult_485_C412_n305,
         dp_cluster_0_mult_485_C412_n304, dp_cluster_0_mult_485_C412_n303,
         dp_cluster_0_mult_485_C412_n302, dp_cluster_0_mult_485_C412_n301,
         dp_cluster_0_mult_485_C412_n300, dp_cluster_0_mult_485_C412_n299,
         dp_cluster_0_mult_485_C412_n298, dp_cluster_0_mult_485_C412_n297,
         dp_cluster_0_mult_485_C412_n296, dp_cluster_0_mult_485_C412_n295,
         dp_cluster_0_mult_485_C412_n294, dp_cluster_0_mult_485_C412_n293,
         dp_cluster_0_mult_485_C412_n292, dp_cluster_0_mult_485_C412_n291,
         dp_cluster_0_mult_485_C412_n290, dp_cluster_0_mult_485_C412_n289,
         dp_cluster_0_mult_485_C412_n288, dp_cluster_0_mult_485_C412_n287,
         dp_cluster_0_mult_485_C412_n286, dp_cluster_0_mult_485_C412_n285,
         dp_cluster_0_mult_485_C412_n284, dp_cluster_0_mult_485_C412_n283,
         dp_cluster_0_mult_485_C412_n282, dp_cluster_0_mult_485_C412_n281,
         dp_cluster_0_mult_485_C412_n280, dp_cluster_0_mult_485_C412_n279,
         dp_cluster_0_mult_485_C412_n278, dp_cluster_0_mult_485_C412_n277,
         dp_cluster_0_mult_485_C412_n275, dp_cluster_0_mult_485_C412_n274,
         dp_cluster_0_mult_485_C412_n273, dp_cluster_0_mult_485_C412_n272,
         dp_cluster_0_mult_485_C412_n271, dp_cluster_0_mult_485_C412_n270,
         dp_cluster_0_mult_485_C412_n269, dp_cluster_0_mult_485_C412_n268,
         dp_cluster_0_mult_485_C412_n267, dp_cluster_0_mult_485_C412_n266,
         dp_cluster_0_mult_485_C412_n264, dp_cluster_0_mult_485_C412_n263,
         dp_cluster_0_mult_485_C412_n262, dp_cluster_0_mult_485_C412_n261,
         dp_cluster_0_mult_485_C412_n260, dp_cluster_0_mult_485_C412_n259,
         dp_cluster_0_mult_485_C412_n258, dp_cluster_0_mult_485_C412_n257,
         dp_cluster_0_mult_485_C412_n256, dp_cluster_0_mult_485_C412_n255,
         dp_cluster_0_mult_485_C412_n254, dp_cluster_0_mult_485_C412_n253,
         dp_cluster_0_mult_485_C412_n252, dp_cluster_0_mult_485_C412_n250,
         dp_cluster_0_mult_485_C412_n249, dp_cluster_0_mult_485_C412_n248,
         dp_cluster_0_mult_485_C412_n247, dp_cluster_0_mult_485_C412_n246,
         dp_cluster_0_mult_485_C412_n245, dp_cluster_0_mult_485_C412_n244,
         dp_cluster_0_mult_485_C412_n243, dp_cluster_0_mult_485_C412_n242,
         dp_cluster_0_mult_485_C412_n241, dp_cluster_0_mult_485_C412_n240,
         dp_cluster_0_mult_485_C412_n239, dp_cluster_0_mult_485_C412_n238,
         dp_cluster_0_mult_485_C412_n237, dp_cluster_0_mult_485_C412_n236,
         dp_cluster_0_mult_485_C412_n235, dp_cluster_0_mult_485_C412_n234,
         dp_cluster_0_mult_485_C412_n233, dp_cluster_0_mult_485_C412_n232,
         dp_cluster_0_mult_485_C412_n231, dp_cluster_0_mult_485_C412_n230,
         dp_cluster_0_mult_485_C412_n229, dp_cluster_0_mult_485_C412_n228,
         dp_cluster_0_mult_485_C412_n227, dp_cluster_0_mult_485_C412_n226,
         dp_cluster_0_mult_485_C412_n225, dp_cluster_0_mult_485_C412_n224,
         dp_cluster_0_mult_485_C412_n223, dp_cluster_0_mult_485_C412_n222,
         dp_cluster_0_mult_485_C412_n221, dp_cluster_0_mult_485_C412_n220,
         dp_cluster_0_mult_485_C412_n219, dp_cluster_0_mult_485_C412_n218,
         dp_cluster_0_mult_485_C412_n217, dp_cluster_0_mult_485_C412_n216,
         dp_cluster_0_mult_485_C412_n215, dp_cluster_0_mult_485_C412_n214,
         dp_cluster_0_mult_485_C412_n213, dp_cluster_0_mult_485_C412_n212,
         dp_cluster_0_mult_485_C412_n211, dp_cluster_0_mult_485_C412_n210,
         dp_cluster_0_mult_485_C412_n209, dp_cluster_0_mult_485_C412_n208,
         dp_cluster_0_mult_485_C412_n207, dp_cluster_0_mult_485_C412_n206,
         dp_cluster_0_mult_485_C412_n205, dp_cluster_0_mult_485_C412_n204,
         dp_cluster_0_mult_485_C412_n203, dp_cluster_0_mult_485_C412_n202,
         dp_cluster_0_mult_485_C412_n201, dp_cluster_0_mult_485_C412_n200,
         dp_cluster_0_mult_485_C412_n199, dp_cluster_0_mult_485_C412_n198,
         dp_cluster_0_mult_485_C412_n197, dp_cluster_0_mult_485_C412_n196,
         dp_cluster_0_mult_485_C412_n195, dp_cluster_0_mult_485_C412_n194,
         dp_cluster_0_mult_485_C412_n193, dp_cluster_0_mult_485_C412_n192,
         dp_cluster_0_mult_485_C412_n191, dp_cluster_0_mult_485_C412_n190,
         dp_cluster_0_mult_485_C412_n189, dp_cluster_0_mult_485_C412_n188,
         dp_cluster_0_mult_485_C412_n187, dp_cluster_0_mult_485_C412_n186,
         dp_cluster_0_mult_485_C412_n185, dp_cluster_0_mult_485_C412_n184,
         dp_cluster_0_mult_485_C412_n183, dp_cluster_0_mult_485_C412_n182,
         dp_cluster_0_mult_485_C412_n181, dp_cluster_0_mult_485_C412_n180,
         dp_cluster_0_mult_485_C412_n179, dp_cluster_0_mult_485_C412_n178,
         dp_cluster_0_mult_485_C412_n177, dp_cluster_0_mult_485_C412_n176,
         dp_cluster_0_mult_485_C412_n175, dp_cluster_0_mult_485_C412_n174,
         dp_cluster_0_mult_485_C412_n173, dp_cluster_0_mult_485_C412_n172,
         dp_cluster_0_mult_485_C412_n171, dp_cluster_0_mult_485_C412_n170,
         dp_cluster_0_mult_485_C412_n169, dp_cluster_0_mult_485_C412_n168,
         dp_cluster_0_mult_485_C412_n167, dp_cluster_0_mult_485_C412_n166,
         dp_cluster_0_mult_485_C412_n165, dp_cluster_0_mult_485_C412_n164,
         dp_cluster_0_mult_485_C412_n163, dp_cluster_0_mult_485_C412_n162,
         dp_cluster_0_mult_485_C412_n161, dp_cluster_0_mult_485_C412_n160,
         dp_cluster_0_mult_485_C412_n159, dp_cluster_0_mult_485_C412_n158,
         dp_cluster_0_mult_485_C412_n157, dp_cluster_0_mult_485_C412_n156,
         dp_cluster_0_mult_485_C412_n155, dp_cluster_0_mult_485_C412_n154,
         dp_cluster_0_mult_485_C412_n153, dp_cluster_0_mult_485_C412_n152,
         dp_cluster_0_mult_485_C412_n150, dp_cluster_0_mult_485_C412_n149,
         dp_cluster_0_mult_485_C412_n148, dp_cluster_0_mult_485_C412_n147,
         dp_cluster_0_mult_485_C412_n146, dp_cluster_0_mult_485_C412_n145,
         dp_cluster_0_mult_485_C412_n144, dp_cluster_0_mult_485_C412_n143,
         dp_cluster_0_mult_485_C412_n142, dp_cluster_0_mult_485_C412_n141,
         dp_cluster_0_mult_485_C412_n140, dp_cluster_0_mult_485_C412_n139,
         dp_cluster_0_mult_485_C412_n138, dp_cluster_0_mult_485_C412_n137,
         dp_cluster_0_mult_485_C412_n136, dp_cluster_0_mult_485_C412_n135,
         dp_cluster_0_mult_485_C412_n134, dp_cluster_0_mult_485_C412_n133,
         dp_cluster_0_mult_485_C412_n132, dp_cluster_0_mult_485_C412_n130,
         dp_cluster_0_mult_485_C412_n129, dp_cluster_0_mult_485_C412_n128,
         dp_cluster_0_mult_485_C412_n127, dp_cluster_0_mult_485_C412_n126,
         dp_cluster_0_mult_485_C412_n125, dp_cluster_0_mult_485_C412_n124,
         dp_cluster_0_mult_485_C412_n123, dp_cluster_0_mult_485_C412_n122,
         dp_cluster_0_mult_485_C412_n121, dp_cluster_0_mult_485_C412_n120,
         dp_cluster_0_mult_485_C412_n119, dp_cluster_0_mult_485_C412_n118,
         dp_cluster_0_mult_485_C412_n117, dp_cluster_0_mult_485_C412_n116,
         dp_cluster_0_mult_485_C412_n115, dp_cluster_0_mult_485_C412_n114,
         dp_cluster_0_mult_485_C412_n112, dp_cluster_0_mult_485_C412_n111,
         dp_cluster_0_mult_485_C412_n110, dp_cluster_0_mult_485_C412_n109,
         dp_cluster_0_mult_485_C412_n108, dp_cluster_0_mult_485_C412_n107,
         dp_cluster_0_mult_485_C412_n106, dp_cluster_0_mult_485_C412_n105,
         dp_cluster_0_mult_485_C412_n104, dp_cluster_0_mult_485_C412_n103,
         dp_cluster_0_mult_485_C412_n102, dp_cluster_0_mult_485_C412_n101,
         dp_cluster_0_mult_485_C412_n100, dp_cluster_0_mult_485_C412_n98,
         dp_cluster_0_mult_485_C412_n97, dp_cluster_0_mult_485_C412_n96,
         dp_cluster_0_mult_485_C412_n95, dp_cluster_0_mult_485_C412_n94,
         dp_cluster_0_mult_485_C412_n93, dp_cluster_0_mult_485_C412_n92,
         dp_cluster_0_mult_485_C412_n91, dp_cluster_0_mult_485_C412_n90,
         dp_cluster_0_mult_485_C412_n89, dp_cluster_0_mult_485_C412_n88,
         dp_cluster_0_mult_485_C412_n86, dp_cluster_0_mult_485_C412_n85,
         dp_cluster_0_mult_485_C412_n84, dp_cluster_0_mult_485_C412_n83,
         dp_cluster_0_mult_485_C412_n82, dp_cluster_0_mult_485_C412_n81,
         dp_cluster_0_mult_485_C412_n80, dp_cluster_0_mult_485_C412_n77,
         dp_cluster_0_mult_485_C412_n76, dp_cluster_0_mult_485_C412_n75,
         dp_cluster_0_mult_485_C412_n74, dp_cluster_0_mult_485_C412_n73,
         dp_cluster_0_mult_485_C412_n72, dp_cluster_0_mult_485_C412_n71,
         dp_cluster_0_mult_485_C412_n70, dp_cluster_0_mult_485_C412_n69,
         dp_cluster_0_mult_485_C412_n68, dp_cluster_0_mult_485_C412_n67,
         dp_cluster_0_mult_485_C412_n66, dp_cluster_0_mult_485_C412_n65,
         dp_cluster_0_mult_485_C412_n64, dp_cluster_0_mult_485_C412_n63,
         dp_cluster_0_mult_485_C412_n62, dp_cluster_0_mult_485_C412_n61,
         dp_cluster_0_mult_485_C412_n60, dp_cluster_0_mult_485_C412_n59,
         dp_cluster_0_mult_485_C412_n58, dp_cluster_0_mult_485_C412_n57,
         dp_cluster_0_mult_485_C412_n56, dp_cluster_0_mult_485_C412_n55,
         dp_cluster_0_mult_485_C412_n54, dp_cluster_0_mult_485_C412_n53,
         dp_cluster_0_mult_485_C412_n52, dp_cluster_0_mult_486_C412_n376,
         dp_cluster_0_mult_486_C412_n375, dp_cluster_0_mult_486_C412_n374,
         dp_cluster_0_mult_486_C412_n373, dp_cluster_0_mult_486_C412_n372,
         dp_cluster_0_mult_486_C412_n371, dp_cluster_0_mult_486_C412_n370,
         dp_cluster_0_mult_486_C412_n369, dp_cluster_0_mult_486_C412_n368,
         dp_cluster_0_mult_486_C412_n367, dp_cluster_0_mult_486_C412_n366,
         dp_cluster_0_mult_486_C412_n365, dp_cluster_0_mult_486_C412_n364,
         dp_cluster_0_mult_486_C412_n363, dp_cluster_0_mult_486_C412_n362,
         dp_cluster_0_mult_486_C412_n361, dp_cluster_0_mult_486_C412_n360,
         dp_cluster_0_mult_486_C412_n359, dp_cluster_0_mult_486_C412_n358,
         dp_cluster_0_mult_486_C412_n357, dp_cluster_0_mult_486_C412_n356,
         dp_cluster_0_mult_486_C412_n355, dp_cluster_0_mult_486_C412_n354,
         dp_cluster_0_mult_486_C412_n353, dp_cluster_0_mult_486_C412_n352,
         dp_cluster_0_mult_486_C412_n351, dp_cluster_0_mult_486_C412_n350,
         dp_cluster_0_mult_486_C412_n349, dp_cluster_0_mult_486_C412_n348,
         dp_cluster_0_mult_486_C412_n347, dp_cluster_0_mult_486_C412_n346,
         dp_cluster_0_mult_486_C412_n345, dp_cluster_0_mult_486_C412_n344,
         dp_cluster_0_mult_486_C412_n343, dp_cluster_0_mult_486_C412_n342,
         dp_cluster_0_mult_486_C412_n341, dp_cluster_0_mult_486_C412_n340,
         dp_cluster_0_mult_486_C412_n339, dp_cluster_0_mult_486_C412_n338,
         dp_cluster_0_mult_486_C412_n337, dp_cluster_0_mult_486_C412_n336,
         dp_cluster_0_mult_486_C412_n335, dp_cluster_0_mult_486_C412_n334,
         dp_cluster_0_mult_486_C412_n333, dp_cluster_0_mult_486_C412_n332,
         dp_cluster_0_mult_486_C412_n331, dp_cluster_0_mult_486_C412_n330,
         dp_cluster_0_mult_486_C412_n329, dp_cluster_0_mult_486_C412_n328,
         dp_cluster_0_mult_486_C412_n327, dp_cluster_0_mult_486_C412_n326,
         dp_cluster_0_mult_486_C412_n325, dp_cluster_0_mult_486_C412_n324,
         dp_cluster_0_mult_486_C412_n323, dp_cluster_0_mult_486_C412_n322,
         dp_cluster_0_mult_486_C412_n321, dp_cluster_0_mult_486_C412_n320,
         dp_cluster_0_mult_486_C412_n319, dp_cluster_0_mult_486_C412_n317,
         dp_cluster_0_mult_486_C412_n316, dp_cluster_0_mult_486_C412_n315,
         dp_cluster_0_mult_486_C412_n314, dp_cluster_0_mult_486_C412_n313,
         dp_cluster_0_mult_486_C412_n312, dp_cluster_0_mult_486_C412_n311,
         dp_cluster_0_mult_486_C412_n310, dp_cluster_0_mult_486_C412_n309,
         dp_cluster_0_mult_486_C412_n308, dp_cluster_0_mult_486_C412_n307,
         dp_cluster_0_mult_486_C412_n306, dp_cluster_0_mult_486_C412_n305,
         dp_cluster_0_mult_486_C412_n304, dp_cluster_0_mult_486_C412_n303,
         dp_cluster_0_mult_486_C412_n302, dp_cluster_0_mult_486_C412_n301,
         dp_cluster_0_mult_486_C412_n300, dp_cluster_0_mult_486_C412_n299,
         dp_cluster_0_mult_486_C412_n298, dp_cluster_0_mult_486_C412_n297,
         dp_cluster_0_mult_486_C412_n296, dp_cluster_0_mult_486_C412_n295,
         dp_cluster_0_mult_486_C412_n294, dp_cluster_0_mult_486_C412_n293,
         dp_cluster_0_mult_486_C412_n292, dp_cluster_0_mult_486_C412_n291,
         dp_cluster_0_mult_486_C412_n290, dp_cluster_0_mult_486_C412_n289,
         dp_cluster_0_mult_486_C412_n288, dp_cluster_0_mult_486_C412_n287,
         dp_cluster_0_mult_486_C412_n286, dp_cluster_0_mult_486_C412_n285,
         dp_cluster_0_mult_486_C412_n284, dp_cluster_0_mult_486_C412_n283,
         dp_cluster_0_mult_486_C412_n282, dp_cluster_0_mult_486_C412_n281,
         dp_cluster_0_mult_486_C412_n280, dp_cluster_0_mult_486_C412_n279,
         dp_cluster_0_mult_486_C412_n278, dp_cluster_0_mult_486_C412_n277,
         dp_cluster_0_mult_486_C412_n275, dp_cluster_0_mult_486_C412_n274,
         dp_cluster_0_mult_486_C412_n273, dp_cluster_0_mult_486_C412_n272,
         dp_cluster_0_mult_486_C412_n271, dp_cluster_0_mult_486_C412_n270,
         dp_cluster_0_mult_486_C412_n269, dp_cluster_0_mult_486_C412_n268,
         dp_cluster_0_mult_486_C412_n267, dp_cluster_0_mult_486_C412_n266,
         dp_cluster_0_mult_486_C412_n264, dp_cluster_0_mult_486_C412_n263,
         dp_cluster_0_mult_486_C412_n262, dp_cluster_0_mult_486_C412_n261,
         dp_cluster_0_mult_486_C412_n260, dp_cluster_0_mult_486_C412_n259,
         dp_cluster_0_mult_486_C412_n258, dp_cluster_0_mult_486_C412_n257,
         dp_cluster_0_mult_486_C412_n256, dp_cluster_0_mult_486_C412_n255,
         dp_cluster_0_mult_486_C412_n254, dp_cluster_0_mult_486_C412_n253,
         dp_cluster_0_mult_486_C412_n252, dp_cluster_0_mult_486_C412_n250,
         dp_cluster_0_mult_486_C412_n249, dp_cluster_0_mult_486_C412_n248,
         dp_cluster_0_mult_486_C412_n247, dp_cluster_0_mult_486_C412_n246,
         dp_cluster_0_mult_486_C412_n245, dp_cluster_0_mult_486_C412_n244,
         dp_cluster_0_mult_486_C412_n243, dp_cluster_0_mult_486_C412_n242,
         dp_cluster_0_mult_486_C412_n241, dp_cluster_0_mult_486_C412_n240,
         dp_cluster_0_mult_486_C412_n239, dp_cluster_0_mult_486_C412_n238,
         dp_cluster_0_mult_486_C412_n237, dp_cluster_0_mult_486_C412_n236,
         dp_cluster_0_mult_486_C412_n235, dp_cluster_0_mult_486_C412_n234,
         dp_cluster_0_mult_486_C412_n233, dp_cluster_0_mult_486_C412_n232,
         dp_cluster_0_mult_486_C412_n231, dp_cluster_0_mult_486_C412_n230,
         dp_cluster_0_mult_486_C412_n229, dp_cluster_0_mult_486_C412_n228,
         dp_cluster_0_mult_486_C412_n227, dp_cluster_0_mult_486_C412_n226,
         dp_cluster_0_mult_486_C412_n225, dp_cluster_0_mult_486_C412_n224,
         dp_cluster_0_mult_486_C412_n223, dp_cluster_0_mult_486_C412_n222,
         dp_cluster_0_mult_486_C412_n221, dp_cluster_0_mult_486_C412_n220,
         dp_cluster_0_mult_486_C412_n219, dp_cluster_0_mult_486_C412_n218,
         dp_cluster_0_mult_486_C412_n217, dp_cluster_0_mult_486_C412_n216,
         dp_cluster_0_mult_486_C412_n215, dp_cluster_0_mult_486_C412_n214,
         dp_cluster_0_mult_486_C412_n213, dp_cluster_0_mult_486_C412_n212,
         dp_cluster_0_mult_486_C412_n211, dp_cluster_0_mult_486_C412_n210,
         dp_cluster_0_mult_486_C412_n209, dp_cluster_0_mult_486_C412_n208,
         dp_cluster_0_mult_486_C412_n207, dp_cluster_0_mult_486_C412_n206,
         dp_cluster_0_mult_486_C412_n205, dp_cluster_0_mult_486_C412_n204,
         dp_cluster_0_mult_486_C412_n203, dp_cluster_0_mult_486_C412_n202,
         dp_cluster_0_mult_486_C412_n201, dp_cluster_0_mult_486_C412_n200,
         dp_cluster_0_mult_486_C412_n199, dp_cluster_0_mult_486_C412_n198,
         dp_cluster_0_mult_486_C412_n197, dp_cluster_0_mult_486_C412_n196,
         dp_cluster_0_mult_486_C412_n195, dp_cluster_0_mult_486_C412_n194,
         dp_cluster_0_mult_486_C412_n193, dp_cluster_0_mult_486_C412_n192,
         dp_cluster_0_mult_486_C412_n191, dp_cluster_0_mult_486_C412_n190,
         dp_cluster_0_mult_486_C412_n189, dp_cluster_0_mult_486_C412_n188,
         dp_cluster_0_mult_486_C412_n187, dp_cluster_0_mult_486_C412_n186,
         dp_cluster_0_mult_486_C412_n185, dp_cluster_0_mult_486_C412_n184,
         dp_cluster_0_mult_486_C412_n183, dp_cluster_0_mult_486_C412_n182,
         dp_cluster_0_mult_486_C412_n181, dp_cluster_0_mult_486_C412_n180,
         dp_cluster_0_mult_486_C412_n179, dp_cluster_0_mult_486_C412_n178,
         dp_cluster_0_mult_486_C412_n177, dp_cluster_0_mult_486_C412_n176,
         dp_cluster_0_mult_486_C412_n175, dp_cluster_0_mult_486_C412_n174,
         dp_cluster_0_mult_486_C412_n173, dp_cluster_0_mult_486_C412_n172,
         dp_cluster_0_mult_486_C412_n171, dp_cluster_0_mult_486_C412_n170,
         dp_cluster_0_mult_486_C412_n169, dp_cluster_0_mult_486_C412_n168,
         dp_cluster_0_mult_486_C412_n167, dp_cluster_0_mult_486_C412_n166,
         dp_cluster_0_mult_486_C412_n165, dp_cluster_0_mult_486_C412_n164,
         dp_cluster_0_mult_486_C412_n163, dp_cluster_0_mult_486_C412_n162,
         dp_cluster_0_mult_486_C412_n161, dp_cluster_0_mult_486_C412_n160,
         dp_cluster_0_mult_486_C412_n159, dp_cluster_0_mult_486_C412_n158,
         dp_cluster_0_mult_486_C412_n157, dp_cluster_0_mult_486_C412_n156,
         dp_cluster_0_mult_486_C412_n155, dp_cluster_0_mult_486_C412_n154,
         dp_cluster_0_mult_486_C412_n153, dp_cluster_0_mult_486_C412_n152,
         dp_cluster_0_mult_486_C412_n150, dp_cluster_0_mult_486_C412_n149,
         dp_cluster_0_mult_486_C412_n148, dp_cluster_0_mult_486_C412_n147,
         dp_cluster_0_mult_486_C412_n146, dp_cluster_0_mult_486_C412_n145,
         dp_cluster_0_mult_486_C412_n144, dp_cluster_0_mult_486_C412_n143,
         dp_cluster_0_mult_486_C412_n142, dp_cluster_0_mult_486_C412_n141,
         dp_cluster_0_mult_486_C412_n140, dp_cluster_0_mult_486_C412_n139,
         dp_cluster_0_mult_486_C412_n138, dp_cluster_0_mult_486_C412_n137,
         dp_cluster_0_mult_486_C412_n136, dp_cluster_0_mult_486_C412_n135,
         dp_cluster_0_mult_486_C412_n134, dp_cluster_0_mult_486_C412_n133,
         dp_cluster_0_mult_486_C412_n132, dp_cluster_0_mult_486_C412_n130,
         dp_cluster_0_mult_486_C412_n129, dp_cluster_0_mult_486_C412_n128,
         dp_cluster_0_mult_486_C412_n127, dp_cluster_0_mult_486_C412_n126,
         dp_cluster_0_mult_486_C412_n125, dp_cluster_0_mult_486_C412_n124,
         dp_cluster_0_mult_486_C412_n123, dp_cluster_0_mult_486_C412_n122,
         dp_cluster_0_mult_486_C412_n121, dp_cluster_0_mult_486_C412_n120,
         dp_cluster_0_mult_486_C412_n119, dp_cluster_0_mult_486_C412_n118,
         dp_cluster_0_mult_486_C412_n117, dp_cluster_0_mult_486_C412_n116,
         dp_cluster_0_mult_486_C412_n115, dp_cluster_0_mult_486_C412_n114,
         dp_cluster_0_mult_486_C412_n112, dp_cluster_0_mult_486_C412_n111,
         dp_cluster_0_mult_486_C412_n110, dp_cluster_0_mult_486_C412_n109,
         dp_cluster_0_mult_486_C412_n108, dp_cluster_0_mult_486_C412_n107,
         dp_cluster_0_mult_486_C412_n106, dp_cluster_0_mult_486_C412_n105,
         dp_cluster_0_mult_486_C412_n104, dp_cluster_0_mult_486_C412_n103,
         dp_cluster_0_mult_486_C412_n102, dp_cluster_0_mult_486_C412_n101,
         dp_cluster_0_mult_486_C412_n100, dp_cluster_0_mult_486_C412_n98,
         dp_cluster_0_mult_486_C412_n97, dp_cluster_0_mult_486_C412_n96,
         dp_cluster_0_mult_486_C412_n95, dp_cluster_0_mult_486_C412_n94,
         dp_cluster_0_mult_486_C412_n93, dp_cluster_0_mult_486_C412_n92,
         dp_cluster_0_mult_486_C412_n91, dp_cluster_0_mult_486_C412_n90,
         dp_cluster_0_mult_486_C412_n89, dp_cluster_0_mult_486_C412_n88,
         dp_cluster_0_mult_486_C412_n86, dp_cluster_0_mult_486_C412_n85,
         dp_cluster_0_mult_486_C412_n84, dp_cluster_0_mult_486_C412_n83,
         dp_cluster_0_mult_486_C412_n82, dp_cluster_0_mult_486_C412_n81,
         dp_cluster_0_mult_486_C412_n80, dp_cluster_0_mult_486_C412_n77,
         dp_cluster_0_mult_486_C412_n76, dp_cluster_0_mult_486_C412_n75,
         dp_cluster_0_mult_486_C412_n74, dp_cluster_0_mult_486_C412_n73,
         dp_cluster_0_mult_486_C412_n72, dp_cluster_0_mult_486_C412_n71,
         dp_cluster_0_mult_486_C412_n70, dp_cluster_0_mult_486_C412_n69,
         dp_cluster_0_mult_486_C412_n68, dp_cluster_0_mult_486_C412_n67,
         dp_cluster_0_mult_486_C412_n66, dp_cluster_0_mult_486_C412_n65,
         dp_cluster_0_mult_486_C412_n64, dp_cluster_0_mult_486_C412_n63,
         dp_cluster_0_mult_486_C412_n62, dp_cluster_0_mult_486_C412_n61,
         dp_cluster_0_mult_486_C412_n60, dp_cluster_0_mult_486_C412_n59,
         dp_cluster_0_mult_486_C412_n58, dp_cluster_0_mult_486_C412_n57,
         dp_cluster_0_mult_486_C412_n56, dp_cluster_0_mult_486_C412_n55,
         dp_cluster_0_mult_486_C412_n54, dp_cluster_0_mult_486_C412_n53,
         dp_cluster_0_mult_486_C412_n52, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987;
  wire   [15:0] xo0_r_w_d1r;
  wire   [15:0] xo0_i_w_d1r;
  wire   [15:0] xo1_r_w_d1r;
  wire   [15:0] xo1_i_w_d1r;
  wire   [15:0] xo2_r_w_d1r;
  wire   [15:0] xo2_i_w_d1r;
  wire   [15:0] xo3_r_w_d1r;
  wire   [15:0] xo3_i_w_d1r;
  wire   [15:0] xo4_r_w_d1r;
  wire   [15:0] xo4_i_w_d1r;
  wire   [15:0] xo5_r_w_d1r;
  wire   [15:0] xo5_i_w_d1r;
  wire   [15:0] xo6_r_w_d1r;
  wire   [15:0] xo6_i_w_d1r;
  wire   [15:0] xo7_r_w_d1r;
  wire   [15:0] xo7_i_w_d1r;
  wire   [16:1] s1_0_r;
  wire   [16:1] s1_0_i;
  wire   [16:1] s1_1_r;
  wire   [16:1] s1_1_i;
  wire   [16:1] s1_2_r;
  wire   [16:1] s1_2_i;
  wire   [16:1] s1_3_r;
  wire   [16:1] s1_3_i;
  wire   [15:0] s1_5_tmp_r;
  wire   [15:0] s1_5_tmp_i;
  wire   [15:0] s1_6_tmp_i;
  wire   [15:0] s1_7_tmp_r;
  wire   [15:0] s1_7_tmp_i;
  wire   [16:1] s1_4_r;
  wire   [16:1] s1_5_r;
  wire   [16:2] s1_6_r;
  wire   [16:1] s1_7_r;
  wire   [16:1] s1_4_i;
  wire   [16:1] s1_5_i;
  wire   [16:1] s1_6_i;
  wire   [16:1] s1_7_i;
  wire   [15:0] s2_0_r;
  wire   [15:0] s2_1_r;
  wire   [15:0] s2_2_r;
  wire   [15:0] s2_4_r;
  wire   [15:0] s2_5_r;
  wire   [15:0] s2_6_r;
  wire   [15:0] s2_0_i;
  wire   [15:0] s2_1_i;
  wire   [15:0] s2_2_i;
  wire   [15:0] s2_3_i;
  wire   [15:0] s2_4_i;
  wire   [15:0] s2_5_i;
  wire   [15:0] s2_6_i;
  wire   [15:0] s2_7_i;
  wire   [15:0] s3_0_r;
  wire   [15:0] s3_1_r;
  wire   [15:0] s3_2_r;
  wire   [15:0] s3_3_r;
  wire   [15:0] s3_4_r;
  wire   [15:0] s3_5_r;
  wire   [15:0] s3_6_r;
  wire   [15:0] s3_7_r;
  wire   [15:0] s3_0_i;
  wire   [15:0] s3_1_i;
  wire   [15:0] s3_2_i;
  wire   [15:0] s3_3_i;
  wire   [15:0] s3_4_i;
  wire   [15:0] s3_5_i;
  wire   [15:0] s3_6_i;
  wire   [15:0] s3_7_i;
  wire   [15:1] dp_cluster_4_s2_7_r;
  wire   [15:1] dp_cluster_5_s2_3_r;
  wire   [15:1] dp_cluster_5_sub_1_root_sub_440_carry;
  wire   [15:1] dp_cluster_4_sub_1_root_sub_444_carry;
  wire   [27:12] dp_cluster_3_add_514_C415_carry;
  wire   [27:12] dp_cluster_2_sub_487_C409_carry;
  wire   [27:12] dp_cluster_1_add_514_C418_carry;
  wire   [27:12] dp_cluster_0_sub_487_C412_carry;
  wire   [15:1] sub_385_carry;
  wire   [15:2] add_384_carry;
  wire   [15:1] sub_383_carry;
  wire   [15:2] add_382_carry;
  wire   [15:1] sub_381_carry;
  wire   [15:2] add_380_carry;
  wire   [15:1] sub_379_carry;
  wire   [15:2] add_378_carry;
  wire   [15:1] sub_376_carry;
  wire   [15:2] add_375_carry;
  wire   [15:1] sub_374_carry;
  wire   [15:2] add_373_carry;
  wire   [15:1] sub_372_carry;
  wire   [15:2] add_371_carry;
  wire   [15:1] sub_370_carry;
  wire   [15:2] add_369_carry;
  wire   [15:1] sub_365_carry;
  wire   [15:1] sub_364_carry;
  wire   [15:2] add_363_carry;
  wire   [15:2] add_362_carry;
  wire   [15:1] sub_361_carry;
  wire   [15:1] sub_360_carry;
  wire   [15:2] add_359_carry;
  wire   [15:2] add_358_carry;
  wire   [15:1] sub_355_carry;
  wire   [15:2] add_354_carry;
  wire   [15:2] add_353_carry;
  wire   [15:1] sub_351_carry;
  wire   [15:2] add_350_carry;
  wire   [15:2] add_349_carry;
  wire   [16:1] sub_344_carry;
  wire   [16:1] sub_343_carry;
  wire   [16:1] sub_342_carry;
  wire   [16:1] sub_341_carry;
  wire   [16:1] add_340_carry;
  wire   [16:1] add_339_carry;
  wire   [16:1] add_338_carry;
  wire   [16:1] add_337_carry;
  wire   [16:1] sub_335_carry;
  wire   [16:1] sub_334_carry;
  wire   [16:1] sub_333_carry;
  wire   [16:1] sub_332_carry;
  wire   [16:1] add_331_carry;
  wire   [16:1] add_330_carry;
  wire   [16:1] add_329_carry;
  wire   [16:1] add_328_carry;

  DFCNQD1 valid_in_d1r_reg ( .D(valid_in), .CP(clk), .CDN(reset_n), .Q(
        valid_in_d1r) );
  DFCNQD1 valid_in_d2r_reg ( .D(valid_in_d1r), .CP(clk), .CDN(reset_n), .Q(
        valid_out) );
  DFCNQD1 xo0_r_w_d1r_reg_15_ ( .D(s1_0_r[16]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[15]) );
  DFCNQD1 xo0_r_w_d1r_reg_14_ ( .D(s1_0_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[14]) );
  DFCNQD1 xo0_r_w_d1r_reg_13_ ( .D(s1_0_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[13]) );
  DFCNQD1 xo0_r_w_d1r_reg_12_ ( .D(s1_0_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[12]) );
  DFCNQD1 xo0_r_w_d1r_reg_11_ ( .D(s1_0_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[11]) );
  DFCNQD1 xo0_r_w_d1r_reg_10_ ( .D(s1_0_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[10]) );
  DFCNQD1 xo0_r_w_d1r_reg_9_ ( .D(s1_0_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[9]) );
  DFCNQD1 xo0_r_w_d1r_reg_8_ ( .D(s1_0_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[8]) );
  DFCNQD1 xo0_r_w_d1r_reg_7_ ( .D(s1_0_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[7]) );
  DFCNQD1 xo0_r_w_d1r_reg_6_ ( .D(s1_0_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[6]) );
  DFCNQD1 xo0_r_w_d1r_reg_5_ ( .D(s1_0_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[5]) );
  DFCNQD1 xo0_r_w_d1r_reg_4_ ( .D(s1_0_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[4]) );
  DFCNQD1 xo0_r_w_d1r_reg_3_ ( .D(s1_0_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[3]) );
  DFCNQD1 xo0_r_w_d1r_reg_2_ ( .D(s1_0_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[2]) );
  DFCNQD1 xo0_r_w_d1r_reg_1_ ( .D(s1_0_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[1]) );
  DFCNQD1 xo0_r_w_d1r_reg_0_ ( .D(s1_0_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r_w_d1r[0]) );
  DFCNQD1 xo0_i_w_d1r_reg_15_ ( .D(s1_0_i[16]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[15]) );
  DFCNQD1 xo0_i_w_d1r_reg_14_ ( .D(s1_0_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[14]) );
  DFCNQD1 xo0_i_w_d1r_reg_13_ ( .D(s1_0_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[13]) );
  DFCNQD1 xo0_i_w_d1r_reg_12_ ( .D(s1_0_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[12]) );
  DFCNQD1 xo0_i_w_d1r_reg_11_ ( .D(s1_0_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[11]) );
  DFCNQD1 xo0_i_w_d1r_reg_10_ ( .D(s1_0_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[10]) );
  DFCNQD1 xo0_i_w_d1r_reg_9_ ( .D(s1_0_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[9]) );
  DFCNQD1 xo0_i_w_d1r_reg_8_ ( .D(s1_0_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[8]) );
  DFCNQD1 xo0_i_w_d1r_reg_7_ ( .D(s1_0_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[7]) );
  DFCNQD1 xo0_i_w_d1r_reg_6_ ( .D(s1_0_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[6]) );
  DFCNQD1 xo0_i_w_d1r_reg_5_ ( .D(s1_0_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[5]) );
  DFCNQD1 xo0_i_w_d1r_reg_4_ ( .D(s1_0_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[4]) );
  DFCNQD1 xo0_i_w_d1r_reg_3_ ( .D(s1_0_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[3]) );
  DFCNQD1 xo0_i_w_d1r_reg_2_ ( .D(s1_0_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[2]) );
  DFCNQD1 xo0_i_w_d1r_reg_1_ ( .D(s1_0_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[1]) );
  DFCNQD1 xo0_i_w_d1r_reg_0_ ( .D(s1_0_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i_w_d1r[0]) );
  DFCNQD1 xo1_r_w_d1r_reg_15_ ( .D(s1_1_r[16]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[15]) );
  DFCNQD1 xo1_r_w_d1r_reg_14_ ( .D(s1_1_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[14]) );
  DFCNQD1 xo1_r_w_d1r_reg_13_ ( .D(s1_1_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[13]) );
  DFCNQD1 xo1_r_w_d1r_reg_12_ ( .D(s1_1_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[12]) );
  DFCNQD1 xo1_r_w_d1r_reg_11_ ( .D(s1_1_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[11]) );
  DFCNQD1 xo1_r_w_d1r_reg_10_ ( .D(s1_1_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[10]) );
  DFCNQD1 xo1_r_w_d1r_reg_9_ ( .D(s1_1_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[9]) );
  DFCNQD1 xo1_r_w_d1r_reg_8_ ( .D(s1_1_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[8]) );
  DFCNQD1 xo1_r_w_d1r_reg_7_ ( .D(s1_1_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[7]) );
  DFCNQD1 xo1_r_w_d1r_reg_6_ ( .D(s1_1_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[6]) );
  DFCNQD1 xo1_r_w_d1r_reg_5_ ( .D(s1_1_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[5]) );
  DFCNQD1 xo1_r_w_d1r_reg_4_ ( .D(s1_1_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[4]) );
  DFCNQD1 xo1_r_w_d1r_reg_3_ ( .D(s1_1_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[3]) );
  DFCNQD1 xo1_r_w_d1r_reg_2_ ( .D(s1_1_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[2]) );
  DFCNQD1 xo1_r_w_d1r_reg_1_ ( .D(s1_1_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[1]) );
  DFCNQD1 xo1_r_w_d1r_reg_0_ ( .D(s1_1_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r_w_d1r[0]) );
  DFCNQD1 xo1_i_w_d1r_reg_15_ ( .D(s1_1_i[16]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[15]) );
  DFCNQD1 xo1_i_w_d1r_reg_14_ ( .D(s1_1_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[14]) );
  DFCNQD1 xo1_i_w_d1r_reg_13_ ( .D(s1_1_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[13]) );
  DFCNQD1 xo1_i_w_d1r_reg_12_ ( .D(s1_1_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[12]) );
  DFCNQD1 xo1_i_w_d1r_reg_11_ ( .D(s1_1_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[11]) );
  DFCNQD1 xo1_i_w_d1r_reg_10_ ( .D(s1_1_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[10]) );
  DFCNQD1 xo1_i_w_d1r_reg_9_ ( .D(s1_1_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[9]) );
  DFCNQD1 xo1_i_w_d1r_reg_8_ ( .D(s1_1_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[8]) );
  DFCNQD1 xo1_i_w_d1r_reg_7_ ( .D(s1_1_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[7]) );
  DFCNQD1 xo1_i_w_d1r_reg_6_ ( .D(s1_1_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[6]) );
  DFCNQD1 xo1_i_w_d1r_reg_5_ ( .D(s1_1_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[5]) );
  DFCNQD1 xo1_i_w_d1r_reg_4_ ( .D(s1_1_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[4]) );
  DFCNQD1 xo1_i_w_d1r_reg_3_ ( .D(s1_1_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[3]) );
  DFCNQD1 xo1_i_w_d1r_reg_2_ ( .D(s1_1_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[2]) );
  DFCNQD1 xo1_i_w_d1r_reg_1_ ( .D(s1_1_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[1]) );
  DFCNQD1 xo1_i_w_d1r_reg_0_ ( .D(s1_1_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i_w_d1r[0]) );
  DFCNQD1 xo2_r_w_d1r_reg_15_ ( .D(s1_2_r[16]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[15]) );
  DFCNQD1 xo2_r_w_d1r_reg_14_ ( .D(s1_2_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[14]) );
  DFCNQD1 xo2_r_w_d1r_reg_13_ ( .D(s1_2_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[13]) );
  DFCNQD1 xo2_r_w_d1r_reg_12_ ( .D(s1_2_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[12]) );
  DFCNQD1 xo2_r_w_d1r_reg_11_ ( .D(s1_2_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[11]) );
  DFCNQD1 xo2_r_w_d1r_reg_10_ ( .D(s1_2_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[10]) );
  DFCNQD1 xo2_r_w_d1r_reg_9_ ( .D(s1_2_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[9]) );
  DFCNQD1 xo2_r_w_d1r_reg_8_ ( .D(s1_2_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[8]) );
  DFCNQD1 xo2_r_w_d1r_reg_7_ ( .D(s1_2_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[7]) );
  DFCNQD1 xo2_r_w_d1r_reg_6_ ( .D(s1_2_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[6]) );
  DFCNQD1 xo2_r_w_d1r_reg_5_ ( .D(s1_2_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[5]) );
  DFCNQD1 xo2_r_w_d1r_reg_4_ ( .D(s1_2_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[4]) );
  DFCNQD1 xo2_r_w_d1r_reg_3_ ( .D(s1_2_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[3]) );
  DFCNQD1 xo2_r_w_d1r_reg_2_ ( .D(s1_2_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[2]) );
  DFCNQD1 xo2_r_w_d1r_reg_1_ ( .D(s1_2_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[1]) );
  DFCNQD1 xo2_r_w_d1r_reg_0_ ( .D(s1_2_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r_w_d1r[0]) );
  DFCNQD1 xo2_i_w_d1r_reg_15_ ( .D(s1_2_i[16]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[15]) );
  DFCNQD1 xo2_i_w_d1r_reg_14_ ( .D(s1_2_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[14]) );
  DFCNQD1 xo2_i_w_d1r_reg_13_ ( .D(s1_2_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[13]) );
  DFCNQD1 xo2_i_w_d1r_reg_12_ ( .D(s1_2_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[12]) );
  DFCNQD1 xo2_i_w_d1r_reg_11_ ( .D(s1_2_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[11]) );
  DFCNQD1 xo2_i_w_d1r_reg_10_ ( .D(s1_2_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[10]) );
  DFCNQD1 xo2_i_w_d1r_reg_9_ ( .D(s1_2_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[9]) );
  DFCNQD1 xo2_i_w_d1r_reg_8_ ( .D(s1_2_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[8]) );
  DFCNQD1 xo2_i_w_d1r_reg_7_ ( .D(s1_2_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[7]) );
  DFCNQD1 xo2_i_w_d1r_reg_6_ ( .D(s1_2_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[6]) );
  DFCNQD1 xo2_i_w_d1r_reg_5_ ( .D(s1_2_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[5]) );
  DFCNQD1 xo2_i_w_d1r_reg_4_ ( .D(s1_2_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[4]) );
  DFCNQD1 xo2_i_w_d1r_reg_3_ ( .D(s1_2_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[3]) );
  DFCNQD1 xo2_i_w_d1r_reg_2_ ( .D(s1_2_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[2]) );
  DFCNQD1 xo2_i_w_d1r_reg_1_ ( .D(s1_2_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[1]) );
  DFCNQD1 xo2_i_w_d1r_reg_0_ ( .D(s1_2_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i_w_d1r[0]) );
  DFCNQD1 xo3_r_w_d1r_reg_15_ ( .D(s1_3_r[16]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[15]) );
  DFCNQD1 xo3_r_w_d1r_reg_14_ ( .D(s1_3_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[14]) );
  DFCNQD1 xo3_r_w_d1r_reg_13_ ( .D(s1_3_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[13]) );
  DFCNQD1 xo3_r_w_d1r_reg_12_ ( .D(s1_3_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[12]) );
  DFCNQD1 xo3_r_w_d1r_reg_11_ ( .D(s1_3_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[11]) );
  DFCNQD1 xo3_r_w_d1r_reg_10_ ( .D(s1_3_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[10]) );
  DFCNQD1 xo3_r_w_d1r_reg_9_ ( .D(s1_3_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[9]) );
  DFCNQD1 xo3_r_w_d1r_reg_8_ ( .D(s1_3_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[8]) );
  DFCNQD1 xo3_r_w_d1r_reg_7_ ( .D(s1_3_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[7]) );
  DFCNQD1 xo3_r_w_d1r_reg_6_ ( .D(s1_3_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[6]) );
  DFCNQD1 xo3_r_w_d1r_reg_5_ ( .D(s1_3_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[5]) );
  DFCNQD1 xo3_r_w_d1r_reg_4_ ( .D(s1_3_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[4]) );
  DFCNQD1 xo3_r_w_d1r_reg_3_ ( .D(s1_3_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[3]) );
  DFCNQD1 xo3_r_w_d1r_reg_2_ ( .D(s1_3_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[2]) );
  DFCNQD1 xo3_r_w_d1r_reg_1_ ( .D(s1_3_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[1]) );
  DFCNQD1 xo3_r_w_d1r_reg_0_ ( .D(s1_3_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r_w_d1r[0]) );
  DFCNQD1 xo3_i_w_d1r_reg_15_ ( .D(s1_3_i[16]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[15]) );
  DFCNQD1 xo3_i_w_d1r_reg_14_ ( .D(s1_3_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[14]) );
  DFCNQD1 xo3_i_w_d1r_reg_13_ ( .D(s1_3_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[13]) );
  DFCNQD1 xo3_i_w_d1r_reg_12_ ( .D(s1_3_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[12]) );
  DFCNQD1 xo3_i_w_d1r_reg_11_ ( .D(s1_3_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[11]) );
  DFCNQD1 xo3_i_w_d1r_reg_10_ ( .D(s1_3_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[10]) );
  DFCNQD1 xo3_i_w_d1r_reg_9_ ( .D(s1_3_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[9]) );
  DFCNQD1 xo3_i_w_d1r_reg_8_ ( .D(s1_3_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[8]) );
  DFCNQD1 xo3_i_w_d1r_reg_7_ ( .D(s1_3_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[7]) );
  DFCNQD1 xo3_i_w_d1r_reg_6_ ( .D(s1_3_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[6]) );
  DFCNQD1 xo3_i_w_d1r_reg_5_ ( .D(s1_3_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[5]) );
  DFCNQD1 xo3_i_w_d1r_reg_4_ ( .D(s1_3_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[4]) );
  DFCNQD1 xo3_i_w_d1r_reg_3_ ( .D(s1_3_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[3]) );
  DFCNQD1 xo3_i_w_d1r_reg_2_ ( .D(s1_3_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[2]) );
  DFCNQD1 xo3_i_w_d1r_reg_1_ ( .D(s1_3_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[1]) );
  DFCNQD1 xo3_i_w_d1r_reg_0_ ( .D(s1_3_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i_w_d1r[0]) );
  DFCNQD1 xo4_r_w_d1r_reg_15_ ( .D(s1_4_r[16]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[15]) );
  DFCNQD1 xo4_r_w_d1r_reg_14_ ( .D(s1_4_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[14]) );
  DFCNQD1 xo4_r_w_d1r_reg_13_ ( .D(s1_4_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[13]) );
  DFCNQD1 xo4_r_w_d1r_reg_12_ ( .D(s1_4_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[12]) );
  DFCNQD1 xo4_r_w_d1r_reg_11_ ( .D(s1_4_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[11]) );
  DFCNQD1 xo4_r_w_d1r_reg_10_ ( .D(s1_4_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[10]) );
  DFCNQD1 xo4_r_w_d1r_reg_9_ ( .D(s1_4_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[9]) );
  DFCNQD1 xo4_r_w_d1r_reg_8_ ( .D(s1_4_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[8]) );
  DFCNQD1 xo4_r_w_d1r_reg_7_ ( .D(s1_4_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[7]) );
  DFCNQD1 xo4_r_w_d1r_reg_6_ ( .D(s1_4_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[6]) );
  DFCNQD1 xo4_r_w_d1r_reg_5_ ( .D(s1_4_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[5]) );
  DFCNQD1 xo4_r_w_d1r_reg_4_ ( .D(s1_4_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[4]) );
  DFCNQD1 xo4_r_w_d1r_reg_3_ ( .D(s1_4_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[3]) );
  DFCNQD1 xo4_r_w_d1r_reg_2_ ( .D(s1_4_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[2]) );
  DFCNQD1 xo4_r_w_d1r_reg_1_ ( .D(s1_4_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[1]) );
  DFCNQD1 xo4_r_w_d1r_reg_0_ ( .D(s1_4_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r_w_d1r[0]) );
  DFCNQD1 xo4_i_w_d1r_reg_15_ ( .D(s1_4_i[16]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[15]) );
  DFCNQD1 xo4_i_w_d1r_reg_14_ ( .D(s1_4_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[14]) );
  DFCNQD1 xo4_i_w_d1r_reg_13_ ( .D(s1_4_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[13]) );
  DFCNQD1 xo4_i_w_d1r_reg_12_ ( .D(s1_4_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[12]) );
  DFCNQD1 xo4_i_w_d1r_reg_11_ ( .D(s1_4_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[11]) );
  DFCNQD1 xo4_i_w_d1r_reg_10_ ( .D(s1_4_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[10]) );
  DFCNQD1 xo4_i_w_d1r_reg_9_ ( .D(s1_4_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[9]) );
  DFCNQD1 xo4_i_w_d1r_reg_8_ ( .D(s1_4_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[8]) );
  DFCNQD1 xo4_i_w_d1r_reg_7_ ( .D(s1_4_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[7]) );
  DFCNQD1 xo4_i_w_d1r_reg_6_ ( .D(s1_4_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[6]) );
  DFCNQD1 xo4_i_w_d1r_reg_5_ ( .D(s1_4_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[5]) );
  DFCNQD1 xo4_i_w_d1r_reg_4_ ( .D(s1_4_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[4]) );
  DFCNQD1 xo4_i_w_d1r_reg_3_ ( .D(s1_4_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[3]) );
  DFCNQD1 xo4_i_w_d1r_reg_2_ ( .D(s1_4_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[2]) );
  DFCNQD1 xo4_i_w_d1r_reg_1_ ( .D(s1_4_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[1]) );
  DFCNQD1 xo4_i_w_d1r_reg_0_ ( .D(s1_4_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i_w_d1r[0]) );
  DFCNQD1 xo5_r_w_d1r_reg_15_ ( .D(s1_5_tmp_r[15]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_r_w_d1r[15]) );
  DFCNQD1 xo5_r_w_d1r_reg_14_ ( .D(s1_5_tmp_r[14]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_r_w_d1r[14]) );
  DFCNQD1 xo5_r_w_d1r_reg_13_ ( .D(s1_5_tmp_r[13]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_r_w_d1r[13]) );
  DFCNQD1 xo5_r_w_d1r_reg_12_ ( .D(s1_5_tmp_r[12]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_r_w_d1r[12]) );
  DFCNQD1 xo5_r_w_d1r_reg_11_ ( .D(s1_5_tmp_r[11]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_r_w_d1r[11]) );
  DFCNQD1 xo5_r_w_d1r_reg_10_ ( .D(s1_5_tmp_r[10]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_r_w_d1r[10]) );
  DFCNQD1 xo5_r_w_d1r_reg_9_ ( .D(s1_5_tmp_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[9]) );
  DFCNQD1 xo5_r_w_d1r_reg_8_ ( .D(s1_5_tmp_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[8]) );
  DFCNQD1 xo5_r_w_d1r_reg_7_ ( .D(s1_5_tmp_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[7]) );
  DFCNQD1 xo5_r_w_d1r_reg_6_ ( .D(s1_5_tmp_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[6]) );
  DFCNQD1 xo5_r_w_d1r_reg_5_ ( .D(s1_5_tmp_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[5]) );
  DFCNQD1 xo5_r_w_d1r_reg_4_ ( .D(s1_5_tmp_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[4]) );
  DFCNQD1 xo5_r_w_d1r_reg_3_ ( .D(s1_5_tmp_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[3]) );
  DFCNQD1 xo5_r_w_d1r_reg_2_ ( .D(s1_5_tmp_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[2]) );
  DFCNQD1 xo5_r_w_d1r_reg_1_ ( .D(s1_5_tmp_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[1]) );
  DFCNQD1 xo5_r_w_d1r_reg_0_ ( .D(s1_5_tmp_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r_w_d1r[0]) );
  DFCNQD1 xo5_i_w_d1r_reg_15_ ( .D(s1_5_tmp_i[15]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_i_w_d1r[15]) );
  DFCNQD1 xo5_i_w_d1r_reg_14_ ( .D(s1_5_tmp_i[14]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_i_w_d1r[14]) );
  DFCNQD1 xo5_i_w_d1r_reg_13_ ( .D(s1_5_tmp_i[13]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_i_w_d1r[13]) );
  DFCNQD1 xo5_i_w_d1r_reg_12_ ( .D(s1_5_tmp_i[12]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_i_w_d1r[12]) );
  DFCNQD1 xo5_i_w_d1r_reg_11_ ( .D(s1_5_tmp_i[11]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_i_w_d1r[11]) );
  DFCNQD1 xo5_i_w_d1r_reg_10_ ( .D(s1_5_tmp_i[10]), .CP(clk), .CDN(reset_n), 
        .Q(xo5_i_w_d1r[10]) );
  DFCNQD1 xo5_i_w_d1r_reg_9_ ( .D(s1_5_tmp_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[9]) );
  DFCNQD1 xo5_i_w_d1r_reg_8_ ( .D(s1_5_tmp_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[8]) );
  DFCNQD1 xo5_i_w_d1r_reg_7_ ( .D(s1_5_tmp_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[7]) );
  DFCNQD1 xo5_i_w_d1r_reg_6_ ( .D(s1_5_tmp_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[6]) );
  DFCNQD1 xo5_i_w_d1r_reg_5_ ( .D(s1_5_tmp_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[5]) );
  DFCNQD1 xo5_i_w_d1r_reg_4_ ( .D(s1_5_tmp_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[4]) );
  DFCNQD1 xo5_i_w_d1r_reg_3_ ( .D(s1_5_tmp_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[3]) );
  DFCNQD1 xo5_i_w_d1r_reg_2_ ( .D(s1_5_tmp_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[2]) );
  DFCNQD1 xo5_i_w_d1r_reg_1_ ( .D(s1_5_tmp_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[1]) );
  DFCNQD1 xo5_i_w_d1r_reg_0_ ( .D(s1_5_tmp_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i_w_d1r[0]) );
  DFCNQD1 xo6_r_w_d1r_reg_15_ ( .D(s1_6_i[16]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[15]) );
  DFCNQD1 xo6_r_w_d1r_reg_14_ ( .D(s1_6_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[14]) );
  DFCNQD1 xo6_r_w_d1r_reg_13_ ( .D(s1_6_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[13]) );
  DFCNQD1 xo6_r_w_d1r_reg_12_ ( .D(s1_6_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[12]) );
  DFCNQD1 xo6_r_w_d1r_reg_11_ ( .D(s1_6_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[11]) );
  DFCNQD1 xo6_r_w_d1r_reg_10_ ( .D(s1_6_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[10]) );
  DFCNQD1 xo6_r_w_d1r_reg_9_ ( .D(s1_6_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[9]) );
  DFCNQD1 xo6_r_w_d1r_reg_8_ ( .D(s1_6_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[8]) );
  DFCNQD1 xo6_r_w_d1r_reg_7_ ( .D(s1_6_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[7]) );
  DFCNQD1 xo6_r_w_d1r_reg_6_ ( .D(s1_6_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[6]) );
  DFCNQD1 xo6_r_w_d1r_reg_5_ ( .D(s1_6_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[5]) );
  DFCNQD1 xo6_r_w_d1r_reg_4_ ( .D(s1_6_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[4]) );
  DFCNQD1 xo6_r_w_d1r_reg_3_ ( .D(s1_6_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[3]) );
  DFCNQD1 xo6_r_w_d1r_reg_2_ ( .D(s1_6_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[2]) );
  DFCNQD1 xo6_r_w_d1r_reg_1_ ( .D(s1_6_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[1]) );
  DFCNQD1 xo6_r_w_d1r_reg_0_ ( .D(s1_6_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r_w_d1r[0]) );
  DFCNQD1 xo6_i_w_d1r_reg_15_ ( .D(s1_6_tmp_i[15]), .CP(clk), .CDN(reset_n), 
        .Q(xo6_i_w_d1r[15]) );
  DFCNQD1 xo6_i_w_d1r_reg_14_ ( .D(s1_6_tmp_i[14]), .CP(clk), .CDN(reset_n), 
        .Q(xo6_i_w_d1r[14]) );
  DFCNQD1 xo6_i_w_d1r_reg_13_ ( .D(s1_6_tmp_i[13]), .CP(clk), .CDN(reset_n), 
        .Q(xo6_i_w_d1r[13]) );
  DFCNQD1 xo6_i_w_d1r_reg_12_ ( .D(s1_6_tmp_i[12]), .CP(clk), .CDN(reset_n), 
        .Q(xo6_i_w_d1r[12]) );
  DFCNQD1 xo6_i_w_d1r_reg_11_ ( .D(s1_6_tmp_i[11]), .CP(clk), .CDN(reset_n), 
        .Q(xo6_i_w_d1r[11]) );
  DFCNQD1 xo6_i_w_d1r_reg_10_ ( .D(s1_6_tmp_i[10]), .CP(clk), .CDN(reset_n), 
        .Q(xo6_i_w_d1r[10]) );
  DFCNQD1 xo6_i_w_d1r_reg_9_ ( .D(s1_6_tmp_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[9]) );
  DFCNQD1 xo6_i_w_d1r_reg_8_ ( .D(s1_6_tmp_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[8]) );
  DFCNQD1 xo6_i_w_d1r_reg_7_ ( .D(s1_6_tmp_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[7]) );
  DFCNQD1 xo6_i_w_d1r_reg_6_ ( .D(s1_6_tmp_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[6]) );
  DFCNQD1 xo6_i_w_d1r_reg_5_ ( .D(s1_6_tmp_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[5]) );
  DFCNQD1 xo6_i_w_d1r_reg_4_ ( .D(s1_6_tmp_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[4]) );
  DFCNQD1 xo6_i_w_d1r_reg_3_ ( .D(s1_6_tmp_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[3]) );
  DFCNQD1 xo6_i_w_d1r_reg_2_ ( .D(s1_6_tmp_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[2]) );
  DFCNQD1 xo6_i_w_d1r_reg_1_ ( .D(s1_6_tmp_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[1]) );
  DFCNQD1 xo6_i_w_d1r_reg_0_ ( .D(s1_6_tmp_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i_w_d1r[0]) );
  DFCNQD1 xo7_r_w_d1r_reg_15_ ( .D(s1_7_tmp_r[15]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_r_w_d1r[15]) );
  DFCNQD1 xo7_r_w_d1r_reg_14_ ( .D(s1_7_tmp_r[14]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_r_w_d1r[14]) );
  DFCNQD1 xo7_r_w_d1r_reg_13_ ( .D(s1_7_tmp_r[13]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_r_w_d1r[13]) );
  DFCNQD1 xo7_r_w_d1r_reg_12_ ( .D(s1_7_tmp_r[12]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_r_w_d1r[12]) );
  DFCNQD1 xo7_r_w_d1r_reg_11_ ( .D(s1_7_tmp_r[11]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_r_w_d1r[11]) );
  DFCNQD1 xo7_r_w_d1r_reg_10_ ( .D(s1_7_tmp_r[10]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_r_w_d1r[10]) );
  DFCNQD1 xo7_r_w_d1r_reg_9_ ( .D(s1_7_tmp_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[9]) );
  DFCNQD1 xo7_r_w_d1r_reg_8_ ( .D(s1_7_tmp_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[8]) );
  DFCNQD1 xo7_r_w_d1r_reg_7_ ( .D(s1_7_tmp_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[7]) );
  DFCNQD1 xo7_r_w_d1r_reg_6_ ( .D(s1_7_tmp_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[6]) );
  DFCNQD1 xo7_r_w_d1r_reg_5_ ( .D(s1_7_tmp_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[5]) );
  DFCNQD1 xo7_r_w_d1r_reg_4_ ( .D(s1_7_tmp_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[4]) );
  DFCNQD1 xo7_r_w_d1r_reg_3_ ( .D(s1_7_tmp_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[3]) );
  DFCNQD1 xo7_r_w_d1r_reg_2_ ( .D(s1_7_tmp_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[2]) );
  DFCNQD1 xo7_r_w_d1r_reg_1_ ( .D(s1_7_tmp_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[1]) );
  DFCNQD1 xo7_r_w_d1r_reg_0_ ( .D(s1_7_tmp_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r_w_d1r[0]) );
  DFCNQD1 xo7_i_w_d2r_reg_0_ ( .D(s3_7_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[48]) );
  DFCNQD1 xo7_i_w_d2r_reg_1_ ( .D(s3_7_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[49]) );
  DFCNQD1 xo7_i_w_d2r_reg_2_ ( .D(s3_7_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[50]) );
  DFCNQD1 xo7_i_w_d2r_reg_3_ ( .D(s3_7_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[51]) );
  DFCNQD1 xo7_i_w_d2r_reg_4_ ( .D(s3_7_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[52]) );
  DFCNQD1 xo7_i_w_d2r_reg_5_ ( .D(s3_7_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[53]) );
  DFCNQD1 xo7_i_w_d2r_reg_6_ ( .D(s3_7_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[54]) );
  DFCNQD1 xo7_i_w_d2r_reg_7_ ( .D(s3_7_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[55]) );
  DFCNQD1 xo7_i_w_d2r_reg_8_ ( .D(s3_7_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[56]) );
  DFCNQD1 xo7_i_w_d2r_reg_9_ ( .D(s3_7_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[57]) );
  DFCNQD1 xo7_i_w_d2r_reg_10_ ( .D(s3_7_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[58]) );
  DFCNQD1 xo7_i_w_d2r_reg_11_ ( .D(s3_7_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[59]) );
  DFCNQD1 xo7_i_w_d2r_reg_12_ ( .D(s3_7_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[60]) );
  DFCNQD1 xo7_i_w_d2r_reg_13_ ( .D(s3_7_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[61]) );
  DFCNQD1 xo7_i_w_d2r_reg_14_ ( .D(s3_7_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[62]) );
  DFCNQD1 xo7_i_w_d2r_reg_15_ ( .D(s3_7_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i[63]) );
  DFCNQD1 xo7_i_w_d1r_reg_15_ ( .D(s1_7_tmp_i[15]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_i_w_d1r[15]) );
  DFCNQD1 xo7_i_w_d1r_reg_14_ ( .D(s1_7_tmp_i[14]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_i_w_d1r[14]) );
  DFCNQD1 xo7_i_w_d1r_reg_13_ ( .D(s1_7_tmp_i[13]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_i_w_d1r[13]) );
  DFCNQD1 xo7_i_w_d1r_reg_12_ ( .D(s1_7_tmp_i[12]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_i_w_d1r[12]) );
  DFCNQD1 xo7_i_w_d1r_reg_11_ ( .D(s1_7_tmp_i[11]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_i_w_d1r[11]) );
  DFCNQD1 xo7_i_w_d1r_reg_10_ ( .D(s1_7_tmp_i[10]), .CP(clk), .CDN(reset_n), 
        .Q(xo7_i_w_d1r[10]) );
  DFCNQD1 xo7_i_w_d1r_reg_9_ ( .D(s1_7_tmp_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[9]) );
  DFCNQD1 xo7_i_w_d1r_reg_8_ ( .D(s1_7_tmp_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[8]) );
  DFCNQD1 xo7_i_w_d1r_reg_7_ ( .D(s1_7_tmp_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[7]) );
  DFCNQD1 xo7_i_w_d1r_reg_6_ ( .D(s1_7_tmp_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[6]) );
  DFCNQD1 xo7_i_w_d1r_reg_5_ ( .D(s1_7_tmp_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[5]) );
  DFCNQD1 xo7_i_w_d1r_reg_4_ ( .D(s1_7_tmp_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[4]) );
  DFCNQD1 xo7_i_w_d1r_reg_3_ ( .D(s1_7_tmp_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[3]) );
  DFCNQD1 xo7_i_w_d1r_reg_2_ ( .D(s1_7_tmp_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[2]) );
  DFCNQD1 xo7_i_w_d1r_reg_1_ ( .D(s1_7_tmp_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[1]) );
  DFCNQD1 xo7_i_w_d1r_reg_0_ ( .D(s1_7_tmp_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo7_i_w_d1r[0]) );
  DFCNQD1 xo7_r_w_d2r_reg_0_ ( .D(s3_7_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[48]) );
  DFCNQD1 xo7_r_w_d2r_reg_1_ ( .D(s3_7_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[49]) );
  DFCNQD1 xo7_r_w_d2r_reg_2_ ( .D(s3_7_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[50]) );
  DFCNQD1 xo7_r_w_d2r_reg_3_ ( .D(s3_7_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[51]) );
  DFCNQD1 xo7_r_w_d2r_reg_4_ ( .D(s3_7_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[52]) );
  DFCNQD1 xo7_r_w_d2r_reg_5_ ( .D(s3_7_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[53]) );
  DFCNQD1 xo7_r_w_d2r_reg_6_ ( .D(s3_7_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[54]) );
  DFCNQD1 xo7_r_w_d2r_reg_7_ ( .D(s3_7_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[55]) );
  DFCNQD1 xo7_r_w_d2r_reg_8_ ( .D(s3_7_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[56]) );
  DFCNQD1 xo7_r_w_d2r_reg_9_ ( .D(s3_7_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[57]) );
  DFCNQD1 xo7_r_w_d2r_reg_10_ ( .D(s3_7_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[58]) );
  DFCNQD1 xo7_r_w_d2r_reg_11_ ( .D(s3_7_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[59]) );
  DFCNQD1 xo7_r_w_d2r_reg_12_ ( .D(s3_7_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[60]) );
  DFCNQD1 xo7_r_w_d2r_reg_13_ ( .D(s3_7_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[61]) );
  DFCNQD1 xo7_r_w_d2r_reg_14_ ( .D(s3_7_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[62]) );
  DFCNQD1 xo7_r_w_d2r_reg_15_ ( .D(s3_7_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo7_r[63]) );
  DFCNQD1 xo0_r_w_d2r_reg_15_ ( .D(s3_0_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[63]) );
  DFCNQD1 xo0_r_w_d2r_reg_14_ ( .D(s3_0_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[62]) );
  DFCNQD1 xo0_r_w_d2r_reg_13_ ( .D(s3_0_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[61]) );
  DFCNQD1 xo0_r_w_d2r_reg_12_ ( .D(s3_0_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[60]) );
  DFCNQD1 xo0_r_w_d2r_reg_11_ ( .D(s3_0_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[59]) );
  DFCNQD1 xo0_r_w_d2r_reg_10_ ( .D(s3_0_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[58]) );
  DFCNQD1 xo0_r_w_d2r_reg_9_ ( .D(s3_0_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[57]) );
  DFCNQD1 xo0_r_w_d2r_reg_8_ ( .D(s3_0_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[56]) );
  DFCNQD1 xo0_r_w_d2r_reg_7_ ( .D(s3_0_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[55]) );
  DFCNQD1 xo0_r_w_d2r_reg_6_ ( .D(s3_0_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[54]) );
  DFCNQD1 xo0_r_w_d2r_reg_5_ ( .D(s3_0_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[53]) );
  DFCNQD1 xo0_r_w_d2r_reg_4_ ( .D(s3_0_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[52]) );
  DFCNQD1 xo0_r_w_d2r_reg_3_ ( .D(s3_0_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[51]) );
  DFCNQD1 xo0_r_w_d2r_reg_2_ ( .D(s3_0_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[50]) );
  DFCNQD1 xo0_r_w_d2r_reg_1_ ( .D(s3_0_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[49]) );
  DFCNQD1 xo0_r_w_d2r_reg_0_ ( .D(s3_0_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo0_r[48]) );
  DFCNQD1 xo0_i_w_d2r_reg_15_ ( .D(s3_0_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[63]) );
  DFCNQD1 xo0_i_w_d2r_reg_14_ ( .D(s3_0_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[62]) );
  DFCNQD1 xo0_i_w_d2r_reg_13_ ( .D(s3_0_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[61]) );
  DFCNQD1 xo0_i_w_d2r_reg_12_ ( .D(s3_0_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[60]) );
  DFCNQD1 xo0_i_w_d2r_reg_11_ ( .D(s3_0_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[59]) );
  DFCNQD1 xo0_i_w_d2r_reg_10_ ( .D(s3_0_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[58]) );
  DFCNQD1 xo0_i_w_d2r_reg_9_ ( .D(s3_0_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[57]) );
  DFCNQD1 xo0_i_w_d2r_reg_8_ ( .D(s3_0_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[56]) );
  DFCNQD1 xo0_i_w_d2r_reg_7_ ( .D(s3_0_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[55]) );
  DFCNQD1 xo0_i_w_d2r_reg_6_ ( .D(s3_0_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[54]) );
  DFCNQD1 xo0_i_w_d2r_reg_5_ ( .D(s3_0_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[53]) );
  DFCNQD1 xo0_i_w_d2r_reg_4_ ( .D(s3_0_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[52]) );
  DFCNQD1 xo0_i_w_d2r_reg_3_ ( .D(s3_0_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[51]) );
  DFCNQD1 xo0_i_w_d2r_reg_2_ ( .D(s3_0_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[50]) );
  DFCNQD1 xo0_i_w_d2r_reg_1_ ( .D(s3_0_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[49]) );
  DFCNQD1 xo0_i_w_d2r_reg_0_ ( .D(s3_0_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo0_i[48]) );
  DFCNQD1 xo1_r_w_d2r_reg_15_ ( .D(s3_1_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[63]) );
  DFCNQD1 xo1_r_w_d2r_reg_14_ ( .D(s3_1_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[62]) );
  DFCNQD1 xo1_r_w_d2r_reg_13_ ( .D(s3_1_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[61]) );
  DFCNQD1 xo1_r_w_d2r_reg_12_ ( .D(s3_1_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[60]) );
  DFCNQD1 xo1_r_w_d2r_reg_11_ ( .D(s3_1_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[59]) );
  DFCNQD1 xo1_r_w_d2r_reg_10_ ( .D(s3_1_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[58]) );
  DFCNQD1 xo1_r_w_d2r_reg_9_ ( .D(s3_1_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[57]) );
  DFCNQD1 xo1_r_w_d2r_reg_8_ ( .D(s3_1_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[56]) );
  DFCNQD1 xo1_r_w_d2r_reg_7_ ( .D(s3_1_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[55]) );
  DFCNQD1 xo1_r_w_d2r_reg_6_ ( .D(s3_1_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[54]) );
  DFCNQD1 xo1_r_w_d2r_reg_5_ ( .D(s3_1_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[53]) );
  DFCNQD1 xo1_r_w_d2r_reg_4_ ( .D(s3_1_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[52]) );
  DFCNQD1 xo1_r_w_d2r_reg_3_ ( .D(s3_1_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[51]) );
  DFCNQD1 xo1_r_w_d2r_reg_2_ ( .D(s3_1_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[50]) );
  DFCNQD1 xo1_r_w_d2r_reg_1_ ( .D(s3_1_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[49]) );
  DFCNQD1 xo1_r_w_d2r_reg_0_ ( .D(s3_1_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo1_r[48]) );
  DFCNQD1 xo1_i_w_d2r_reg_15_ ( .D(s3_1_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[63]) );
  DFCNQD1 xo1_i_w_d2r_reg_14_ ( .D(s3_1_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[62]) );
  DFCNQD1 xo1_i_w_d2r_reg_13_ ( .D(s3_1_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[61]) );
  DFCNQD1 xo1_i_w_d2r_reg_12_ ( .D(s3_1_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[60]) );
  DFCNQD1 xo1_i_w_d2r_reg_11_ ( .D(s3_1_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[59]) );
  DFCNQD1 xo1_i_w_d2r_reg_10_ ( .D(s3_1_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[58]) );
  DFCNQD1 xo1_i_w_d2r_reg_9_ ( .D(s3_1_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[57]) );
  DFCNQD1 xo1_i_w_d2r_reg_8_ ( .D(s3_1_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[56]) );
  DFCNQD1 xo1_i_w_d2r_reg_7_ ( .D(s3_1_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[55]) );
  DFCNQD1 xo1_i_w_d2r_reg_6_ ( .D(s3_1_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[54]) );
  DFCNQD1 xo1_i_w_d2r_reg_5_ ( .D(s3_1_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[53]) );
  DFCNQD1 xo1_i_w_d2r_reg_4_ ( .D(s3_1_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[52]) );
  DFCNQD1 xo1_i_w_d2r_reg_3_ ( .D(s3_1_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[51]) );
  DFCNQD1 xo1_i_w_d2r_reg_2_ ( .D(s3_1_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[50]) );
  DFCNQD1 xo1_i_w_d2r_reg_1_ ( .D(s3_1_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[49]) );
  DFCNQD1 xo1_i_w_d2r_reg_0_ ( .D(s3_1_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo1_i[48]) );
  DFCNQD1 xo2_r_w_d2r_reg_15_ ( .D(s3_2_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[63]) );
  DFCNQD1 xo2_r_w_d2r_reg_14_ ( .D(s3_2_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[62]) );
  DFCNQD1 xo2_r_w_d2r_reg_13_ ( .D(s3_2_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[61]) );
  DFCNQD1 xo2_r_w_d2r_reg_12_ ( .D(s3_2_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[60]) );
  DFCNQD1 xo2_r_w_d2r_reg_11_ ( .D(s3_2_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[59]) );
  DFCNQD1 xo2_r_w_d2r_reg_10_ ( .D(s3_2_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[58]) );
  DFCNQD1 xo2_r_w_d2r_reg_9_ ( .D(s3_2_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[57]) );
  DFCNQD1 xo2_r_w_d2r_reg_8_ ( .D(s3_2_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[56]) );
  DFCNQD1 xo2_r_w_d2r_reg_7_ ( .D(s3_2_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[55]) );
  DFCNQD1 xo2_r_w_d2r_reg_6_ ( .D(s3_2_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[54]) );
  DFCNQD1 xo2_r_w_d2r_reg_5_ ( .D(s3_2_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[53]) );
  DFCNQD1 xo2_r_w_d2r_reg_4_ ( .D(s3_2_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[52]) );
  DFCNQD1 xo2_r_w_d2r_reg_3_ ( .D(s3_2_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[51]) );
  DFCNQD1 xo2_r_w_d2r_reg_2_ ( .D(s3_2_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[50]) );
  DFCNQD1 xo2_r_w_d2r_reg_1_ ( .D(s3_2_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[49]) );
  DFCNQD1 xo2_r_w_d2r_reg_0_ ( .D(s3_2_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo2_r[48]) );
  DFCNQD1 xo2_i_w_d2r_reg_15_ ( .D(s3_2_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[63]) );
  DFCNQD1 xo2_i_w_d2r_reg_14_ ( .D(s3_2_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[62]) );
  DFCNQD1 xo2_i_w_d2r_reg_13_ ( .D(s3_2_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[61]) );
  DFCNQD1 xo2_i_w_d2r_reg_12_ ( .D(s3_2_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[60]) );
  DFCNQD1 xo2_i_w_d2r_reg_11_ ( .D(s3_2_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[59]) );
  DFCNQD1 xo2_i_w_d2r_reg_10_ ( .D(s3_2_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[58]) );
  DFCNQD1 xo2_i_w_d2r_reg_9_ ( .D(s3_2_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[57]) );
  DFCNQD1 xo2_i_w_d2r_reg_8_ ( .D(s3_2_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[56]) );
  DFCNQD1 xo2_i_w_d2r_reg_7_ ( .D(s3_2_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[55]) );
  DFCNQD1 xo2_i_w_d2r_reg_6_ ( .D(s3_2_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[54]) );
  DFCNQD1 xo2_i_w_d2r_reg_5_ ( .D(s3_2_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[53]) );
  DFCNQD1 xo2_i_w_d2r_reg_4_ ( .D(s3_2_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[52]) );
  DFCNQD1 xo2_i_w_d2r_reg_3_ ( .D(s3_2_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[51]) );
  DFCNQD1 xo2_i_w_d2r_reg_2_ ( .D(s3_2_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[50]) );
  DFCNQD1 xo2_i_w_d2r_reg_1_ ( .D(s3_2_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[49]) );
  DFCNQD1 xo2_i_w_d2r_reg_0_ ( .D(s3_2_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo2_i[48]) );
  DFCNQD1 xo3_r_w_d2r_reg_15_ ( .D(s3_3_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[63]) );
  DFCNQD1 xo3_r_w_d2r_reg_14_ ( .D(s3_3_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[62]) );
  DFCNQD1 xo3_r_w_d2r_reg_13_ ( .D(s3_3_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[61]) );
  DFCNQD1 xo3_r_w_d2r_reg_12_ ( .D(s3_3_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[60]) );
  DFCNQD1 xo3_r_w_d2r_reg_11_ ( .D(s3_3_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[59]) );
  DFCNQD1 xo3_r_w_d2r_reg_10_ ( .D(s3_3_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[58]) );
  DFCNQD1 xo3_r_w_d2r_reg_9_ ( .D(s3_3_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[57]) );
  DFCNQD1 xo3_r_w_d2r_reg_8_ ( .D(s3_3_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[56]) );
  DFCNQD1 xo3_r_w_d2r_reg_7_ ( .D(s3_3_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[55]) );
  DFCNQD1 xo3_r_w_d2r_reg_6_ ( .D(s3_3_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[54]) );
  DFCNQD1 xo3_r_w_d2r_reg_5_ ( .D(s3_3_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[53]) );
  DFCNQD1 xo3_r_w_d2r_reg_4_ ( .D(s3_3_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[52]) );
  DFCNQD1 xo3_r_w_d2r_reg_3_ ( .D(s3_3_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[51]) );
  DFCNQD1 xo3_r_w_d2r_reg_2_ ( .D(s3_3_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[50]) );
  DFCNQD1 xo3_r_w_d2r_reg_1_ ( .D(s3_3_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[49]) );
  DFCNQD1 xo3_r_w_d2r_reg_0_ ( .D(s3_3_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo3_r[48]) );
  DFCNQD1 xo3_i_w_d2r_reg_15_ ( .D(s3_3_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[63]) );
  DFCNQD1 xo3_i_w_d2r_reg_14_ ( .D(s3_3_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[62]) );
  DFCNQD1 xo3_i_w_d2r_reg_13_ ( .D(s3_3_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[61]) );
  DFCNQD1 xo3_i_w_d2r_reg_12_ ( .D(s3_3_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[60]) );
  DFCNQD1 xo3_i_w_d2r_reg_11_ ( .D(s3_3_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[59]) );
  DFCNQD1 xo3_i_w_d2r_reg_10_ ( .D(s3_3_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[58]) );
  DFCNQD1 xo3_i_w_d2r_reg_9_ ( .D(s3_3_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[57]) );
  DFCNQD1 xo3_i_w_d2r_reg_8_ ( .D(s3_3_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[56]) );
  DFCNQD1 xo3_i_w_d2r_reg_7_ ( .D(s3_3_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[55]) );
  DFCNQD1 xo3_i_w_d2r_reg_6_ ( .D(s3_3_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[54]) );
  DFCNQD1 xo3_i_w_d2r_reg_5_ ( .D(s3_3_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[53]) );
  DFCNQD1 xo3_i_w_d2r_reg_4_ ( .D(s3_3_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[52]) );
  DFCNQD1 xo3_i_w_d2r_reg_3_ ( .D(s3_3_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[51]) );
  DFCNQD1 xo3_i_w_d2r_reg_2_ ( .D(s3_3_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[50]) );
  DFCNQD1 xo3_i_w_d2r_reg_1_ ( .D(s3_3_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[49]) );
  DFCNQD1 xo3_i_w_d2r_reg_0_ ( .D(s3_3_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo3_i[48]) );
  DFCNQD1 xo4_r_w_d2r_reg_15_ ( .D(s3_4_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[63]) );
  DFCNQD1 xo4_r_w_d2r_reg_14_ ( .D(s3_4_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[62]) );
  DFCNQD1 xo4_r_w_d2r_reg_13_ ( .D(s3_4_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[61]) );
  DFCNQD1 xo4_r_w_d2r_reg_12_ ( .D(s3_4_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[60]) );
  DFCNQD1 xo4_r_w_d2r_reg_11_ ( .D(s3_4_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[59]) );
  DFCNQD1 xo4_r_w_d2r_reg_10_ ( .D(s3_4_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[58]) );
  DFCNQD1 xo4_r_w_d2r_reg_9_ ( .D(s3_4_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[57]) );
  DFCNQD1 xo4_r_w_d2r_reg_8_ ( .D(s3_4_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[56]) );
  DFCNQD1 xo4_r_w_d2r_reg_7_ ( .D(s3_4_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[55]) );
  DFCNQD1 xo4_r_w_d2r_reg_6_ ( .D(s3_4_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[54]) );
  DFCNQD1 xo4_r_w_d2r_reg_5_ ( .D(s3_4_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[53]) );
  DFCNQD1 xo4_r_w_d2r_reg_4_ ( .D(s3_4_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[52]) );
  DFCNQD1 xo4_r_w_d2r_reg_3_ ( .D(s3_4_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[51]) );
  DFCNQD1 xo4_r_w_d2r_reg_2_ ( .D(s3_4_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[50]) );
  DFCNQD1 xo4_r_w_d2r_reg_1_ ( .D(s3_4_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[49]) );
  DFCNQD1 xo4_r_w_d2r_reg_0_ ( .D(s3_4_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo4_r[48]) );
  DFCNQD1 xo4_i_w_d2r_reg_15_ ( .D(s3_4_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[63]) );
  DFCNQD1 xo4_i_w_d2r_reg_14_ ( .D(s3_4_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[62]) );
  DFCNQD1 xo4_i_w_d2r_reg_13_ ( .D(s3_4_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[61]) );
  DFCNQD1 xo4_i_w_d2r_reg_12_ ( .D(s3_4_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[60]) );
  DFCNQD1 xo4_i_w_d2r_reg_11_ ( .D(s3_4_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[59]) );
  DFCNQD1 xo4_i_w_d2r_reg_10_ ( .D(s3_4_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[58]) );
  DFCNQD1 xo4_i_w_d2r_reg_9_ ( .D(s3_4_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[57]) );
  DFCNQD1 xo4_i_w_d2r_reg_8_ ( .D(s3_4_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[56]) );
  DFCNQD1 xo4_i_w_d2r_reg_7_ ( .D(s3_4_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[55]) );
  DFCNQD1 xo4_i_w_d2r_reg_6_ ( .D(s3_4_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[54]) );
  DFCNQD1 xo4_i_w_d2r_reg_5_ ( .D(s3_4_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[53]) );
  DFCNQD1 xo4_i_w_d2r_reg_4_ ( .D(s3_4_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[52]) );
  DFCNQD1 xo4_i_w_d2r_reg_3_ ( .D(s3_4_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[51]) );
  DFCNQD1 xo4_i_w_d2r_reg_2_ ( .D(s3_4_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[50]) );
  DFCNQD1 xo4_i_w_d2r_reg_1_ ( .D(s3_4_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[49]) );
  DFCNQD1 xo4_i_w_d2r_reg_0_ ( .D(s3_4_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo4_i[48]) );
  DFCNQD1 xo5_r_w_d2r_reg_15_ ( .D(s3_5_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[63]) );
  DFCNQD1 xo5_r_w_d2r_reg_14_ ( .D(s3_5_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[62]) );
  DFCNQD1 xo5_r_w_d2r_reg_13_ ( .D(s3_5_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[61]) );
  DFCNQD1 xo5_r_w_d2r_reg_12_ ( .D(s3_5_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[60]) );
  DFCNQD1 xo5_r_w_d2r_reg_11_ ( .D(s3_5_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[59]) );
  DFCNQD1 xo5_r_w_d2r_reg_10_ ( .D(s3_5_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[58]) );
  DFCNQD1 xo5_r_w_d2r_reg_9_ ( .D(s3_5_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[57]) );
  DFCNQD1 xo5_r_w_d2r_reg_8_ ( .D(s3_5_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[56]) );
  DFCNQD1 xo5_r_w_d2r_reg_7_ ( .D(s3_5_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[55]) );
  DFCNQD1 xo5_r_w_d2r_reg_6_ ( .D(s3_5_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[54]) );
  DFCNQD1 xo5_r_w_d2r_reg_5_ ( .D(s3_5_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[53]) );
  DFCNQD1 xo5_r_w_d2r_reg_4_ ( .D(s3_5_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[52]) );
  DFCNQD1 xo5_r_w_d2r_reg_3_ ( .D(s3_5_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[51]) );
  DFCNQD1 xo5_r_w_d2r_reg_2_ ( .D(s3_5_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[50]) );
  DFCNQD1 xo5_r_w_d2r_reg_1_ ( .D(s3_5_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[49]) );
  DFCNQD1 xo5_r_w_d2r_reg_0_ ( .D(s3_5_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo5_r[48]) );
  DFCNQD1 xo5_i_w_d2r_reg_15_ ( .D(s3_5_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[63]) );
  DFCNQD1 xo5_i_w_d2r_reg_14_ ( .D(s3_5_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[62]) );
  DFCNQD1 xo5_i_w_d2r_reg_13_ ( .D(s3_5_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[61]) );
  DFCNQD1 xo5_i_w_d2r_reg_12_ ( .D(s3_5_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[60]) );
  DFCNQD1 xo5_i_w_d2r_reg_11_ ( .D(s3_5_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[59]) );
  DFCNQD1 xo5_i_w_d2r_reg_10_ ( .D(s3_5_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[58]) );
  DFCNQD1 xo5_i_w_d2r_reg_9_ ( .D(s3_5_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[57]) );
  DFCNQD1 xo5_i_w_d2r_reg_8_ ( .D(s3_5_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[56]) );
  DFCNQD1 xo5_i_w_d2r_reg_7_ ( .D(s3_5_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[55]) );
  DFCNQD1 xo5_i_w_d2r_reg_6_ ( .D(s3_5_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[54]) );
  DFCNQD1 xo5_i_w_d2r_reg_5_ ( .D(s3_5_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[53]) );
  DFCNQD1 xo5_i_w_d2r_reg_4_ ( .D(s3_5_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[52]) );
  DFCNQD1 xo5_i_w_d2r_reg_3_ ( .D(s3_5_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[51]) );
  DFCNQD1 xo5_i_w_d2r_reg_2_ ( .D(s3_5_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[50]) );
  DFCNQD1 xo5_i_w_d2r_reg_1_ ( .D(s3_5_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[49]) );
  DFCNQD1 xo5_i_w_d2r_reg_0_ ( .D(s3_5_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo5_i[48]) );
  DFCNQD1 xo6_r_w_d2r_reg_15_ ( .D(s3_6_r[15]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[63]) );
  DFCNQD1 xo6_r_w_d2r_reg_14_ ( .D(s3_6_r[14]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[62]) );
  DFCNQD1 xo6_r_w_d2r_reg_13_ ( .D(s3_6_r[13]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[61]) );
  DFCNQD1 xo6_r_w_d2r_reg_12_ ( .D(s3_6_r[12]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[60]) );
  DFCNQD1 xo6_r_w_d2r_reg_11_ ( .D(s3_6_r[11]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[59]) );
  DFCNQD1 xo6_r_w_d2r_reg_10_ ( .D(s3_6_r[10]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[58]) );
  DFCNQD1 xo6_r_w_d2r_reg_9_ ( .D(s3_6_r[9]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[57]) );
  DFCNQD1 xo6_r_w_d2r_reg_8_ ( .D(s3_6_r[8]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[56]) );
  DFCNQD1 xo6_r_w_d2r_reg_7_ ( .D(s3_6_r[7]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[55]) );
  DFCNQD1 xo6_r_w_d2r_reg_6_ ( .D(s3_6_r[6]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[54]) );
  DFCNQD1 xo6_r_w_d2r_reg_5_ ( .D(s3_6_r[5]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[53]) );
  DFCNQD1 xo6_r_w_d2r_reg_4_ ( .D(s3_6_r[4]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[52]) );
  DFCNQD1 xo6_r_w_d2r_reg_3_ ( .D(s3_6_r[3]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[51]) );
  DFCNQD1 xo6_r_w_d2r_reg_2_ ( .D(s3_6_r[2]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[50]) );
  DFCNQD1 xo6_r_w_d2r_reg_1_ ( .D(s3_6_r[1]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[49]) );
  DFCNQD1 xo6_r_w_d2r_reg_0_ ( .D(s3_6_r[0]), .CP(clk), .CDN(reset_n), .Q(
        xo6_r[48]) );
  DFCNQD1 xo6_i_w_d2r_reg_15_ ( .D(s3_6_i[15]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[63]) );
  DFCNQD1 xo6_i_w_d2r_reg_14_ ( .D(s3_6_i[14]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[62]) );
  DFCNQD1 xo6_i_w_d2r_reg_13_ ( .D(s3_6_i[13]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[61]) );
  DFCNQD1 xo6_i_w_d2r_reg_12_ ( .D(s3_6_i[12]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[60]) );
  DFCNQD1 xo6_i_w_d2r_reg_11_ ( .D(s3_6_i[11]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[59]) );
  DFCNQD1 xo6_i_w_d2r_reg_10_ ( .D(s3_6_i[10]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[58]) );
  DFCNQD1 xo6_i_w_d2r_reg_9_ ( .D(s3_6_i[9]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[57]) );
  DFCNQD1 xo6_i_w_d2r_reg_8_ ( .D(s3_6_i[8]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[56]) );
  DFCNQD1 xo6_i_w_d2r_reg_7_ ( .D(s3_6_i[7]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[55]) );
  DFCNQD1 xo6_i_w_d2r_reg_6_ ( .D(s3_6_i[6]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[54]) );
  DFCNQD1 xo6_i_w_d2r_reg_5_ ( .D(s3_6_i[5]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[53]) );
  DFCNQD1 xo6_i_w_d2r_reg_4_ ( .D(s3_6_i[4]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[52]) );
  DFCNQD1 xo6_i_w_d2r_reg_3_ ( .D(s3_6_i[3]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[51]) );
  DFCNQD1 xo6_i_w_d2r_reg_2_ ( .D(s3_6_i[2]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[50]) );
  DFCNQD1 xo6_i_w_d2r_reg_1_ ( .D(s3_6_i[1]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[49]) );
  DFCNQD1 xo6_i_w_d2r_reg_0_ ( .D(s3_6_i[0]), .CP(clk), .CDN(reset_n), .Q(
        xo6_i[48]) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U139 ( .A(
        dp_cluster_3_mult_512_C415_n371), .B(dp_cluster_3_mult_512_C415_n328), 
        .C(dp_cluster_3_mult_512_C415_n342), .CIX(
        dp_cluster_3_mult_512_C415_n237), .D(dp_cluster_3_mult_512_C415_n356), 
        .CO(dp_cluster_3_mult_512_C415_n233), .COX(
        dp_cluster_3_mult_512_C415_n232), .S(dp_cluster_3_mult_512_C415_n234)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U137 ( .A(
        dp_cluster_3_mult_512_C415_n341), .B(dp_cluster_3_mult_512_C415_n370), 
        .C(dp_cluster_3_mult_512_C415_n355), .CIX(
        dp_cluster_3_mult_512_C415_n232), .D(dp_cluster_3_mult_512_C415_n231), 
        .CO(dp_cluster_3_mult_512_C415_n228), .COX(
        dp_cluster_3_mult_512_C415_n227), .S(dp_cluster_3_mult_512_C415_n229)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U135 ( .A(
        dp_cluster_3_mult_512_C415_n354), .B(dp_cluster_3_mult_512_C415_n369), 
        .C(dp_cluster_3_mult_512_C415_n230), .CIX(
        dp_cluster_3_mult_512_C415_n226), .D(dp_cluster_3_mult_512_C415_n227), 
        .CO(dp_cluster_3_mult_512_C415_n223), .COX(
        dp_cluster_3_mult_512_C415_n222), .S(dp_cluster_3_mult_512_C415_n224)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U132 ( .A(
        dp_cluster_3_mult_512_C415_n221), .B(dp_cluster_3_mult_512_C415_n368), 
        .C(dp_cluster_3_mult_512_C415_n225), .CIX(
        dp_cluster_3_mult_512_C415_n222), .D(dp_cluster_3_mult_512_C415_n219), 
        .CO(dp_cluster_3_mult_512_C415_n216), .COX(
        dp_cluster_3_mult_512_C415_n215), .S(dp_cluster_3_mult_512_C415_n217)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U131 ( .A(
        dp_cluster_3_mult_512_C415_n324), .B(dp_cluster_3_mult_512_C415_n295), 
        .C(dp_cluster_3_mult_512_C415_n309), .CIX(
        dp_cluster_3_mult_512_C415_n220), .D(dp_cluster_3_mult_512_C415_n338), 
        .CO(dp_cluster_3_mult_512_C415_n213), .COX(
        dp_cluster_3_mult_512_C415_n212), .S(dp_cluster_3_mult_512_C415_n214)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U130 ( .A(
        dp_cluster_3_mult_512_C415_n352), .B(dp_cluster_3_mult_512_C415_n367), 
        .C(dp_cluster_3_mult_512_C415_n218), .CIX(
        dp_cluster_3_mult_512_C415_n214), .D(dp_cluster_3_mult_512_C415_n215), 
        .CO(dp_cluster_3_mult_512_C415_n210), .COX(
        dp_cluster_3_mult_512_C415_n209), .S(dp_cluster_3_mult_512_C415_n211)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U128 ( .A(
        dp_cluster_3_mult_512_C415_n366), .B(dp_cluster_3_mult_512_C415_n337), 
        .C(dp_cluster_3_mult_512_C415_n351), .CIX(
        dp_cluster_3_mult_512_C415_n212), .D(dp_cluster_3_mult_512_C415_n308), 
        .CO(dp_cluster_3_mult_512_C415_n205), .COX(
        dp_cluster_3_mult_512_C415_n204), .S(dp_cluster_3_mult_512_C415_n206)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U127 ( .A(
        dp_cluster_3_mult_512_C415_n208), .B(dp_cluster_3_mult_512_C415_n323), 
        .C(dp_cluster_3_mult_512_C415_n209), .CIX(
        dp_cluster_3_mult_512_C415_n213), .D(dp_cluster_3_mult_512_C415_n206), 
        .CO(dp_cluster_3_mult_512_C415_n202), .COX(
        dp_cluster_3_mult_512_C415_n201), .S(dp_cluster_3_mult_512_C415_n203)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U125 ( .A(
        dp_cluster_3_mult_512_C415_n322), .B(dp_cluster_3_mult_512_C415_n365), 
        .C(dp_cluster_3_mult_512_C415_n350), .CIX(
        dp_cluster_3_mult_512_C415_n200), .D(dp_cluster_3_mult_512_C415_n207), 
        .CO(dp_cluster_3_mult_512_C415_n197), .COX(
        dp_cluster_3_mult_512_C415_n196), .S(dp_cluster_3_mult_512_C415_n198)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U124 ( .A(
        dp_cluster_3_mult_512_C415_n204), .B(dp_cluster_3_mult_512_C415_n336), 
        .C(dp_cluster_3_mult_512_C415_n198), .CIX(
        dp_cluster_3_mult_512_C415_n201), .D(dp_cluster_3_mult_512_C415_n205), 
        .CO(dp_cluster_3_mult_512_C415_n194), .COX(
        dp_cluster_3_mult_512_C415_n193), .S(dp_cluster_3_mult_512_C415_n195)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U121 ( .A(
        dp_cluster_3_mult_512_C415_n306), .B(dp_cluster_3_mult_512_C415_n349), 
        .C(dp_cluster_3_mult_512_C415_n335), .CIX(
        dp_cluster_3_mult_512_C415_n190), .D(dp_cluster_3_mult_512_C415_n192), 
        .CO(dp_cluster_3_mult_512_C415_n187), .COX(
        dp_cluster_3_mult_512_C415_n186), .S(dp_cluster_3_mult_512_C415_n188)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U120 ( .A(
        dp_cluster_3_mult_512_C415_n199), .B(dp_cluster_3_mult_512_C415_n196), 
        .C(dp_cluster_3_mult_512_C415_n188), .CIX(
        dp_cluster_3_mult_512_C415_n193), .D(dp_cluster_3_mult_512_C415_n197), 
        .CO(dp_cluster_3_mult_512_C415_n184), .COX(
        dp_cluster_3_mult_512_C415_n183), .S(dp_cluster_3_mult_512_C415_n185)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U119 ( .A(
        dp_cluster_3_mult_512_C415_n291), .B(dp_cluster_3_mult_512_C415_n264), 
        .C(dp_cluster_3_mult_512_C415_n278), .CIX(
        dp_cluster_3_mult_512_C415_n191), .D(dp_cluster_3_mult_512_C415_n305), 
        .CO(dp_cluster_3_mult_512_C415_n181), .COX(
        dp_cluster_3_mult_512_C415_n180), .S(dp_cluster_3_mult_512_C415_n182)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U118 ( .A(
        dp_cluster_3_mult_512_C415_n363), .B(dp_cluster_3_mult_512_C415_n334), 
        .C(dp_cluster_3_mult_512_C415_n348), .CIX(
        dp_cluster_3_mult_512_C415_n189), .D(dp_cluster_3_mult_512_C415_n320), 
        .CO(dp_cluster_3_mult_512_C415_n178), .COX(
        dp_cluster_3_mult_512_C415_n177), .S(dp_cluster_3_mult_512_C415_n179)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U117 ( .A(
        dp_cluster_3_mult_512_C415_n182), .B(dp_cluster_3_mult_512_C415_n186), 
        .C(dp_cluster_3_mult_512_C415_n179), .CIX(
        dp_cluster_3_mult_512_C415_n183), .D(dp_cluster_3_mult_512_C415_n187), 
        .CO(dp_cluster_3_mult_512_C415_n175), .COX(
        dp_cluster_3_mult_512_C415_n174), .S(dp_cluster_3_mult_512_C415_n176)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U115 ( .A(
        dp_cluster_3_mult_512_C415_n362), .B(dp_cluster_3_mult_512_C415_n304), 
        .C(dp_cluster_3_mult_512_C415_n347), .CIX(
        dp_cluster_3_mult_512_C415_n180), .D(dp_cluster_3_mult_512_C415_n333), 
        .CO(dp_cluster_3_mult_512_C415_n170), .COX(
        dp_cluster_3_mult_512_C415_n169), .S(dp_cluster_3_mult_512_C415_n171)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U114 ( .A(
        dp_cluster_3_mult_512_C415_n277), .B(dp_cluster_3_mult_512_C415_n319), 
        .C(dp_cluster_3_mult_512_C415_n290), .CIX(
        dp_cluster_3_mult_512_C415_n177), .D(dp_cluster_3_mult_512_C415_n173), 
        .CO(dp_cluster_3_mult_512_C415_n167), .COX(
        dp_cluster_3_mult_512_C415_n166), .S(dp_cluster_3_mult_512_C415_n168)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U113 ( .A(
        dp_cluster_3_mult_512_C415_n168), .B(dp_cluster_3_mult_512_C415_n171), 
        .C(dp_cluster_3_mult_512_C415_n178), .CIX(
        dp_cluster_3_mult_512_C415_n174), .D(dp_cluster_3_mult_512_C415_n181), 
        .CO(dp_cluster_3_mult_512_C415_n164), .COX(
        dp_cluster_3_mult_512_C415_n163), .S(dp_cluster_3_mult_512_C415_n165)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U110 ( .A(
        dp_cluster_3_mult_512_C415_n262), .B(dp_cluster_3_mult_512_C415_n289), 
        .C(dp_cluster_3_mult_512_C415_n361), .CIX(
        dp_cluster_3_mult_512_C415_n169), .D(dp_cluster_3_mult_512_C415_n172), 
        .CO(dp_cluster_3_mult_512_C415_n159), .COX(
        dp_cluster_3_mult_512_C415_n158), .S(dp_cluster_3_mult_512_C415_n160)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U109 ( .A(
        dp_cluster_3_mult_512_C415_n303), .B(dp_cluster_3_mult_512_C415_n346), 
        .C(dp_cluster_3_mult_512_C415_n332), .CIX(
        dp_cluster_3_mult_512_C415_n166), .D(dp_cluster_3_mult_512_C415_n162), 
        .CO(dp_cluster_3_mult_512_C415_n156), .COX(
        dp_cluster_3_mult_512_C415_n155), .S(dp_cluster_3_mult_512_C415_n157)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U108 ( .A(
        dp_cluster_3_mult_512_C415_n170), .B(dp_cluster_3_mult_512_C415_n160), 
        .C(dp_cluster_3_mult_512_C415_n167), .CIX(
        dp_cluster_3_mult_512_C415_n163), .D(dp_cluster_3_mult_512_C415_n157), 
        .CO(dp_cluster_3_mult_512_C415_n153), .COX(
        dp_cluster_3_mult_512_C415_n152), .S(dp_cluster_3_mult_512_C415_n154)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U106 ( .A(
        dp_cluster_3_mult_512_C415_n331), .B(dp_cluster_3_mult_512_C415_n275), 
        .C(n1133), .CIX(dp_cluster_3_mult_512_C415_n158), .D(
        dp_cluster_3_mult_512_C415_n161), .CO(dp_cluster_3_mult_512_C415_n148), 
        .COX(dp_cluster_3_mult_512_C415_n147), .S(
        dp_cluster_3_mult_512_C415_n149) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U105 ( .A(
        dp_cluster_3_mult_512_C415_n317), .B(dp_cluster_3_mult_512_C415_n288), 
        .C(dp_cluster_3_mult_512_C415_n302), .CIX(
        dp_cluster_3_mult_512_C415_n155), .D(dp_cluster_3_mult_512_C415_n261), 
        .CO(dp_cluster_3_mult_512_C415_n145), .COX(
        dp_cluster_3_mult_512_C415_n144), .S(dp_cluster_3_mult_512_C415_n146)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U104 ( .A(
        dp_cluster_3_mult_512_C415_n149), .B(dp_cluster_3_mult_512_C415_n146), 
        .C(dp_cluster_3_mult_512_C415_n156), .CIX(
        dp_cluster_3_mult_512_C415_n152), .D(dp_cluster_3_mult_512_C415_n159), 
        .CO(dp_cluster_3_mult_512_C415_n142), .COX(
        dp_cluster_3_mult_512_C415_n141), .S(dp_cluster_3_mult_512_C415_n143)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U103 ( .A(
        dp_cluster_3_mult_512_C415_n150), .B(dp_cluster_3_mult_512_C415_n260), 
        .C(dp_cluster_3_mult_512_C415_n274), .CIX(
        dp_cluster_3_mult_512_C415_n147), .D(dp_cluster_3_mult_512_C415_n345), 
        .CO(dp_cluster_3_mult_512_C415_n139), .COX(
        dp_cluster_3_mult_512_C415_n138), .S(dp_cluster_3_mult_512_C415_n140)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U102 ( .A(
        dp_cluster_3_mult_512_C415_n330), .B(dp_cluster_3_mult_512_C415_n301), 
        .C(dp_cluster_3_mult_512_C415_n316), .CIX(
        dp_cluster_3_mult_512_C415_n144), .D(dp_cluster_3_mult_512_C415_n287), 
        .CO(dp_cluster_3_mult_512_C415_n136), .COX(
        dp_cluster_3_mult_512_C415_n135), .S(dp_cluster_3_mult_512_C415_n137)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U101 ( .A(
        dp_cluster_3_mult_512_C415_n140), .B(dp_cluster_3_mult_512_C415_n137), 
        .C(dp_cluster_3_mult_512_C415_n145), .CIX(
        dp_cluster_3_mult_512_C415_n141), .D(dp_cluster_3_mult_512_C415_n148), 
        .CO(dp_cluster_3_mult_512_C415_n133), .COX(
        dp_cluster_3_mult_512_C415_n132), .S(dp_cluster_3_mult_512_C415_n134)
         );
  CMPE42D1 dp_cluster_3_mult_512_C415_U98 ( .A(dp_cluster_3_mult_512_C415_n259), .B(dp_cluster_3_mult_512_C415_n300), .C(dp_cluster_3_mult_512_C415_n286), 
        .CIX(dp_cluster_3_mult_512_C415_n129), .D(
        dp_cluster_3_mult_512_C415_n135), .CO(dp_cluster_3_mult_512_C415_n126), 
        .COX(dp_cluster_3_mult_512_C415_n125), .S(
        dp_cluster_3_mult_512_C415_n127) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U97 ( .A(dp_cluster_3_mult_512_C415_n139), .B(dp_cluster_3_mult_512_C415_n138), .C(dp_cluster_3_mult_512_C415_n136), 
        .CIX(dp_cluster_3_mult_512_C415_n132), .D(
        dp_cluster_3_mult_512_C415_n127), .CO(dp_cluster_3_mult_512_C415_n123), 
        .COX(dp_cluster_3_mult_512_C415_n122), .S(
        dp_cluster_3_mult_512_C415_n124) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U95 ( .A(dp_cluster_3_mult_512_C415_n314), .B(dp_cluster_3_mult_512_C415_n285), .C(dp_cluster_3_mult_512_C415_n299), 
        .CIX(dp_cluster_3_mult_512_C415_n121), .D(
        dp_cluster_3_mult_512_C415_n272), .CO(dp_cluster_3_mult_512_C415_n118), 
        .COX(dp_cluster_3_mult_512_C415_n117), .S(
        dp_cluster_3_mult_512_C415_n119) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U94 ( .A(dp_cluster_3_mult_512_C415_n128), .B(dp_cluster_3_mult_512_C415_n125), .C(dp_cluster_3_mult_512_C415_n119), 
        .CIX(dp_cluster_3_mult_512_C415_n122), .D(
        dp_cluster_3_mult_512_C415_n126), .CO(dp_cluster_3_mult_512_C415_n115), 
        .COX(dp_cluster_3_mult_512_C415_n114), .S(
        dp_cluster_3_mult_512_C415_n116) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U92 ( .A(dp_cluster_3_mult_512_C415_n313), .B(dp_cluster_3_mult_512_C415_n271), .C(dp_cluster_3_mult_512_C415_n298), 
        .CIX(dp_cluster_3_mult_512_C415_n120), .D(n1118), .CO(
        dp_cluster_3_mult_512_C415_n110), .COX(dp_cluster_3_mult_512_C415_n109), .S(dp_cluster_3_mult_512_C415_n111) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U91 ( .A(dp_cluster_3_mult_512_C415_n117), .B(dp_cluster_3_mult_512_C415_n257), .C(dp_cluster_3_mult_512_C415_n111), 
        .CIX(dp_cluster_3_mult_512_C415_n114), .D(
        dp_cluster_3_mult_512_C415_n118), .CO(dp_cluster_3_mult_512_C415_n107), 
        .COX(dp_cluster_3_mult_512_C415_n106), .S(
        dp_cluster_3_mult_512_C415_n108) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U90 ( .A(dp_cluster_3_mult_512_C415_n297), .B(dp_cluster_3_mult_512_C415_n256), .C(dp_cluster_3_mult_512_C415_n284), 
        .CIX(dp_cluster_3_mult_512_C415_n109), .D(
        dp_cluster_3_mult_512_C415_n312), .CO(dp_cluster_3_mult_512_C415_n104), 
        .COX(dp_cluster_3_mult_512_C415_n103), .S(
        dp_cluster_3_mult_512_C415_n105) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U89 ( .A(dp_cluster_3_mult_512_C415_n112), .B(dp_cluster_3_mult_512_C415_n270), .C(dp_cluster_3_mult_512_C415_n105), 
        .CIX(dp_cluster_3_mult_512_C415_n106), .D(
        dp_cluster_3_mult_512_C415_n110), .CO(dp_cluster_3_mult_512_C415_n101), 
        .COX(dp_cluster_3_mult_512_C415_n100), .S(
        dp_cluster_3_mult_512_C415_n102) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U86 ( .A(dp_cluster_3_mult_512_C415_n103), .B(dp_cluster_3_mult_512_C415_n283), .C(dp_cluster_3_mult_512_C415_n97), 
        .CIX(dp_cluster_3_mult_512_C415_n100), .D(
        dp_cluster_3_mult_512_C415_n104), .CO(dp_cluster_3_mult_512_C415_n94), 
        .COX(dp_cluster_3_mult_512_C415_n93), .S(
        dp_cluster_3_mult_512_C415_n95) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U84 ( .A(dp_cluster_3_mult_512_C415_n98), 
        .B(dp_cluster_3_mult_512_C415_n282), .C(dp_cluster_3_mult_512_C415_n96), .CIX(dp_cluster_3_mult_512_C415_n93), .D(dp_cluster_3_mult_512_C415_n92), 
        .CO(dp_cluster_3_mult_512_C415_n89), .COX(
        dp_cluster_3_mult_512_C415_n88), .S(dp_cluster_3_mult_512_C415_n90) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U82 ( .A(dp_cluster_3_mult_512_C415_n253), .B(dp_cluster_3_mult_512_C415_n267), .C(n1119), .CIX(
        dp_cluster_3_mult_512_C415_n88), .D(dp_cluster_3_mult_512_C415_n91), 
        .CO(dp_cluster_3_mult_512_C415_n84), .COX(
        dp_cluster_3_mult_512_C415_n83), .S(dp_cluster_3_mult_512_C415_n85) );
  CMPE42D1 dp_cluster_3_mult_512_C415_U81 ( .A(dp_cluster_3_mult_512_C415_n266), .B(dp_cluster_3_mult_512_C415_n86), .C(dp_cluster_3_mult_512_C415_n252), 
        .CIX(dp_cluster_3_mult_512_C415_n83), .D(
        dp_cluster_3_mult_512_C415_n281), .CO(dp_cluster_3_mult_512_C415_n81), 
        .COX(dp_cluster_3_mult_512_C415_n80), .S(
        dp_cluster_3_mult_512_C415_n82) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U139 ( .A(
        dp_cluster_3_mult_513_C415_n371), .B(dp_cluster_3_mult_513_C415_n328), 
        .C(dp_cluster_3_mult_513_C415_n342), .CIX(
        dp_cluster_3_mult_513_C415_n237), .D(dp_cluster_3_mult_513_C415_n356), 
        .CO(dp_cluster_3_mult_513_C415_n233), .COX(
        dp_cluster_3_mult_513_C415_n232), .S(dp_cluster_3_mult_513_C415_n234)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U137 ( .A(
        dp_cluster_3_mult_513_C415_n341), .B(dp_cluster_3_mult_513_C415_n370), 
        .C(dp_cluster_3_mult_513_C415_n355), .CIX(
        dp_cluster_3_mult_513_C415_n232), .D(dp_cluster_3_mult_513_C415_n231), 
        .CO(dp_cluster_3_mult_513_C415_n228), .COX(
        dp_cluster_3_mult_513_C415_n227), .S(dp_cluster_3_mult_513_C415_n229)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U135 ( .A(
        dp_cluster_3_mult_513_C415_n354), .B(dp_cluster_3_mult_513_C415_n369), 
        .C(dp_cluster_3_mult_513_C415_n230), .CIX(
        dp_cluster_3_mult_513_C415_n226), .D(dp_cluster_3_mult_513_C415_n227), 
        .CO(dp_cluster_3_mult_513_C415_n223), .COX(
        dp_cluster_3_mult_513_C415_n222), .S(dp_cluster_3_mult_513_C415_n224)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U132 ( .A(
        dp_cluster_3_mult_513_C415_n221), .B(dp_cluster_3_mult_513_C415_n368), 
        .C(dp_cluster_3_mult_513_C415_n225), .CIX(
        dp_cluster_3_mult_513_C415_n222), .D(dp_cluster_3_mult_513_C415_n219), 
        .CO(dp_cluster_3_mult_513_C415_n216), .COX(
        dp_cluster_3_mult_513_C415_n215), .S(dp_cluster_3_mult_513_C415_n217)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U131 ( .A(
        dp_cluster_3_mult_513_C415_n324), .B(dp_cluster_3_mult_513_C415_n295), 
        .C(dp_cluster_3_mult_513_C415_n309), .CIX(
        dp_cluster_3_mult_513_C415_n220), .D(dp_cluster_3_mult_513_C415_n338), 
        .CO(dp_cluster_3_mult_513_C415_n213), .COX(
        dp_cluster_3_mult_513_C415_n212), .S(dp_cluster_3_mult_513_C415_n214)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U130 ( .A(
        dp_cluster_3_mult_513_C415_n352), .B(dp_cluster_3_mult_513_C415_n367), 
        .C(dp_cluster_3_mult_513_C415_n218), .CIX(
        dp_cluster_3_mult_513_C415_n214), .D(dp_cluster_3_mult_513_C415_n215), 
        .CO(dp_cluster_3_mult_513_C415_n210), .COX(
        dp_cluster_3_mult_513_C415_n209), .S(dp_cluster_3_mult_513_C415_n211)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U128 ( .A(
        dp_cluster_3_mult_513_C415_n366), .B(dp_cluster_3_mult_513_C415_n337), 
        .C(dp_cluster_3_mult_513_C415_n351), .CIX(
        dp_cluster_3_mult_513_C415_n212), .D(dp_cluster_3_mult_513_C415_n308), 
        .CO(dp_cluster_3_mult_513_C415_n205), .COX(
        dp_cluster_3_mult_513_C415_n204), .S(dp_cluster_3_mult_513_C415_n206)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U127 ( .A(
        dp_cluster_3_mult_513_C415_n208), .B(dp_cluster_3_mult_513_C415_n323), 
        .C(dp_cluster_3_mult_513_C415_n209), .CIX(
        dp_cluster_3_mult_513_C415_n213), .D(dp_cluster_3_mult_513_C415_n206), 
        .CO(dp_cluster_3_mult_513_C415_n202), .COX(
        dp_cluster_3_mult_513_C415_n201), .S(dp_cluster_3_mult_513_C415_n203)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U125 ( .A(
        dp_cluster_3_mult_513_C415_n322), .B(dp_cluster_3_mult_513_C415_n365), 
        .C(dp_cluster_3_mult_513_C415_n350), .CIX(
        dp_cluster_3_mult_513_C415_n200), .D(dp_cluster_3_mult_513_C415_n207), 
        .CO(dp_cluster_3_mult_513_C415_n197), .COX(
        dp_cluster_3_mult_513_C415_n196), .S(dp_cluster_3_mult_513_C415_n198)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U124 ( .A(
        dp_cluster_3_mult_513_C415_n204), .B(dp_cluster_3_mult_513_C415_n336), 
        .C(dp_cluster_3_mult_513_C415_n198), .CIX(
        dp_cluster_3_mult_513_C415_n201), .D(dp_cluster_3_mult_513_C415_n205), 
        .CO(dp_cluster_3_mult_513_C415_n194), .COX(
        dp_cluster_3_mult_513_C415_n193), .S(dp_cluster_3_mult_513_C415_n195)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U121 ( .A(
        dp_cluster_3_mult_513_C415_n306), .B(dp_cluster_3_mult_513_C415_n349), 
        .C(dp_cluster_3_mult_513_C415_n335), .CIX(
        dp_cluster_3_mult_513_C415_n190), .D(dp_cluster_3_mult_513_C415_n192), 
        .CO(dp_cluster_3_mult_513_C415_n187), .COX(
        dp_cluster_3_mult_513_C415_n186), .S(dp_cluster_3_mult_513_C415_n188)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U120 ( .A(
        dp_cluster_3_mult_513_C415_n199), .B(dp_cluster_3_mult_513_C415_n196), 
        .C(dp_cluster_3_mult_513_C415_n188), .CIX(
        dp_cluster_3_mult_513_C415_n193), .D(dp_cluster_3_mult_513_C415_n197), 
        .CO(dp_cluster_3_mult_513_C415_n184), .COX(
        dp_cluster_3_mult_513_C415_n183), .S(dp_cluster_3_mult_513_C415_n185)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U119 ( .A(
        dp_cluster_3_mult_513_C415_n291), .B(dp_cluster_3_mult_513_C415_n264), 
        .C(dp_cluster_3_mult_513_C415_n278), .CIX(
        dp_cluster_3_mult_513_C415_n191), .D(dp_cluster_3_mult_513_C415_n305), 
        .CO(dp_cluster_3_mult_513_C415_n181), .COX(
        dp_cluster_3_mult_513_C415_n180), .S(dp_cluster_3_mult_513_C415_n182)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U118 ( .A(
        dp_cluster_3_mult_513_C415_n363), .B(dp_cluster_3_mult_513_C415_n334), 
        .C(dp_cluster_3_mult_513_C415_n348), .CIX(
        dp_cluster_3_mult_513_C415_n189), .D(dp_cluster_3_mult_513_C415_n320), 
        .CO(dp_cluster_3_mult_513_C415_n178), .COX(
        dp_cluster_3_mult_513_C415_n177), .S(dp_cluster_3_mult_513_C415_n179)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U117 ( .A(
        dp_cluster_3_mult_513_C415_n182), .B(dp_cluster_3_mult_513_C415_n186), 
        .C(dp_cluster_3_mult_513_C415_n179), .CIX(
        dp_cluster_3_mult_513_C415_n183), .D(dp_cluster_3_mult_513_C415_n187), 
        .CO(dp_cluster_3_mult_513_C415_n175), .COX(
        dp_cluster_3_mult_513_C415_n174), .S(dp_cluster_3_mult_513_C415_n176)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U115 ( .A(
        dp_cluster_3_mult_513_C415_n362), .B(dp_cluster_3_mult_513_C415_n304), 
        .C(dp_cluster_3_mult_513_C415_n347), .CIX(
        dp_cluster_3_mult_513_C415_n180), .D(dp_cluster_3_mult_513_C415_n333), 
        .CO(dp_cluster_3_mult_513_C415_n170), .COX(
        dp_cluster_3_mult_513_C415_n169), .S(dp_cluster_3_mult_513_C415_n171)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U114 ( .A(
        dp_cluster_3_mult_513_C415_n277), .B(dp_cluster_3_mult_513_C415_n319), 
        .C(dp_cluster_3_mult_513_C415_n290), .CIX(
        dp_cluster_3_mult_513_C415_n177), .D(dp_cluster_3_mult_513_C415_n173), 
        .CO(dp_cluster_3_mult_513_C415_n167), .COX(
        dp_cluster_3_mult_513_C415_n166), .S(dp_cluster_3_mult_513_C415_n168)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U113 ( .A(
        dp_cluster_3_mult_513_C415_n168), .B(dp_cluster_3_mult_513_C415_n171), 
        .C(dp_cluster_3_mult_513_C415_n178), .CIX(
        dp_cluster_3_mult_513_C415_n174), .D(dp_cluster_3_mult_513_C415_n181), 
        .CO(dp_cluster_3_mult_513_C415_n164), .COX(
        dp_cluster_3_mult_513_C415_n163), .S(dp_cluster_3_mult_513_C415_n165)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U110 ( .A(
        dp_cluster_3_mult_513_C415_n262), .B(dp_cluster_3_mult_513_C415_n289), 
        .C(dp_cluster_3_mult_513_C415_n361), .CIX(
        dp_cluster_3_mult_513_C415_n169), .D(dp_cluster_3_mult_513_C415_n172), 
        .CO(dp_cluster_3_mult_513_C415_n159), .COX(
        dp_cluster_3_mult_513_C415_n158), .S(dp_cluster_3_mult_513_C415_n160)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U109 ( .A(
        dp_cluster_3_mult_513_C415_n303), .B(dp_cluster_3_mult_513_C415_n346), 
        .C(dp_cluster_3_mult_513_C415_n332), .CIX(
        dp_cluster_3_mult_513_C415_n166), .D(dp_cluster_3_mult_513_C415_n162), 
        .CO(dp_cluster_3_mult_513_C415_n156), .COX(
        dp_cluster_3_mult_513_C415_n155), .S(dp_cluster_3_mult_513_C415_n157)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U108 ( .A(
        dp_cluster_3_mult_513_C415_n170), .B(dp_cluster_3_mult_513_C415_n160), 
        .C(dp_cluster_3_mult_513_C415_n167), .CIX(
        dp_cluster_3_mult_513_C415_n163), .D(dp_cluster_3_mult_513_C415_n157), 
        .CO(dp_cluster_3_mult_513_C415_n153), .COX(
        dp_cluster_3_mult_513_C415_n152), .S(dp_cluster_3_mult_513_C415_n154)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U106 ( .A(
        dp_cluster_3_mult_513_C415_n331), .B(dp_cluster_3_mult_513_C415_n275), 
        .C(n1270), .CIX(dp_cluster_3_mult_513_C415_n158), .D(
        dp_cluster_3_mult_513_C415_n161), .CO(dp_cluster_3_mult_513_C415_n148), 
        .COX(dp_cluster_3_mult_513_C415_n147), .S(
        dp_cluster_3_mult_513_C415_n149) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U105 ( .A(
        dp_cluster_3_mult_513_C415_n317), .B(dp_cluster_3_mult_513_C415_n288), 
        .C(dp_cluster_3_mult_513_C415_n302), .CIX(
        dp_cluster_3_mult_513_C415_n155), .D(dp_cluster_3_mult_513_C415_n261), 
        .CO(dp_cluster_3_mult_513_C415_n145), .COX(
        dp_cluster_3_mult_513_C415_n144), .S(dp_cluster_3_mult_513_C415_n146)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U104 ( .A(
        dp_cluster_3_mult_513_C415_n149), .B(dp_cluster_3_mult_513_C415_n146), 
        .C(dp_cluster_3_mult_513_C415_n156), .CIX(
        dp_cluster_3_mult_513_C415_n152), .D(dp_cluster_3_mult_513_C415_n159), 
        .CO(dp_cluster_3_mult_513_C415_n142), .COX(
        dp_cluster_3_mult_513_C415_n141), .S(dp_cluster_3_mult_513_C415_n143)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U103 ( .A(
        dp_cluster_3_mult_513_C415_n150), .B(dp_cluster_3_mult_513_C415_n260), 
        .C(dp_cluster_3_mult_513_C415_n274), .CIX(
        dp_cluster_3_mult_513_C415_n147), .D(dp_cluster_3_mult_513_C415_n345), 
        .CO(dp_cluster_3_mult_513_C415_n139), .COX(
        dp_cluster_3_mult_513_C415_n138), .S(dp_cluster_3_mult_513_C415_n140)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U102 ( .A(
        dp_cluster_3_mult_513_C415_n330), .B(dp_cluster_3_mult_513_C415_n301), 
        .C(dp_cluster_3_mult_513_C415_n316), .CIX(
        dp_cluster_3_mult_513_C415_n144), .D(dp_cluster_3_mult_513_C415_n287), 
        .CO(dp_cluster_3_mult_513_C415_n136), .COX(
        dp_cluster_3_mult_513_C415_n135), .S(dp_cluster_3_mult_513_C415_n137)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U101 ( .A(
        dp_cluster_3_mult_513_C415_n140), .B(dp_cluster_3_mult_513_C415_n137), 
        .C(dp_cluster_3_mult_513_C415_n145), .CIX(
        dp_cluster_3_mult_513_C415_n141), .D(dp_cluster_3_mult_513_C415_n148), 
        .CO(dp_cluster_3_mult_513_C415_n133), .COX(
        dp_cluster_3_mult_513_C415_n132), .S(dp_cluster_3_mult_513_C415_n134)
         );
  CMPE42D1 dp_cluster_3_mult_513_C415_U98 ( .A(dp_cluster_3_mult_513_C415_n259), .B(dp_cluster_3_mult_513_C415_n300), .C(dp_cluster_3_mult_513_C415_n286), 
        .CIX(dp_cluster_3_mult_513_C415_n129), .D(
        dp_cluster_3_mult_513_C415_n135), .CO(dp_cluster_3_mult_513_C415_n126), 
        .COX(dp_cluster_3_mult_513_C415_n125), .S(
        dp_cluster_3_mult_513_C415_n127) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U97 ( .A(dp_cluster_3_mult_513_C415_n139), .B(dp_cluster_3_mult_513_C415_n138), .C(dp_cluster_3_mult_513_C415_n136), 
        .CIX(dp_cluster_3_mult_513_C415_n132), .D(
        dp_cluster_3_mult_513_C415_n127), .CO(dp_cluster_3_mult_513_C415_n123), 
        .COX(dp_cluster_3_mult_513_C415_n122), .S(
        dp_cluster_3_mult_513_C415_n124) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U95 ( .A(dp_cluster_3_mult_513_C415_n314), .B(dp_cluster_3_mult_513_C415_n285), .C(dp_cluster_3_mult_513_C415_n299), 
        .CIX(dp_cluster_3_mult_513_C415_n121), .D(
        dp_cluster_3_mult_513_C415_n272), .CO(dp_cluster_3_mult_513_C415_n118), 
        .COX(dp_cluster_3_mult_513_C415_n117), .S(
        dp_cluster_3_mult_513_C415_n119) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U94 ( .A(dp_cluster_3_mult_513_C415_n128), .B(dp_cluster_3_mult_513_C415_n125), .C(dp_cluster_3_mult_513_C415_n119), 
        .CIX(dp_cluster_3_mult_513_C415_n122), .D(
        dp_cluster_3_mult_513_C415_n126), .CO(dp_cluster_3_mult_513_C415_n115), 
        .COX(dp_cluster_3_mult_513_C415_n114), .S(
        dp_cluster_3_mult_513_C415_n116) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U92 ( .A(dp_cluster_3_mult_513_C415_n313), .B(dp_cluster_3_mult_513_C415_n271), .C(dp_cluster_3_mult_513_C415_n298), 
        .CIX(dp_cluster_3_mult_513_C415_n120), .D(n1259), .CO(
        dp_cluster_3_mult_513_C415_n110), .COX(dp_cluster_3_mult_513_C415_n109), .S(dp_cluster_3_mult_513_C415_n111) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U91 ( .A(dp_cluster_3_mult_513_C415_n117), .B(dp_cluster_3_mult_513_C415_n257), .C(dp_cluster_3_mult_513_C415_n111), 
        .CIX(dp_cluster_3_mult_513_C415_n114), .D(
        dp_cluster_3_mult_513_C415_n118), .CO(dp_cluster_3_mult_513_C415_n107), 
        .COX(dp_cluster_3_mult_513_C415_n106), .S(
        dp_cluster_3_mult_513_C415_n108) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U90 ( .A(dp_cluster_3_mult_513_C415_n297), .B(dp_cluster_3_mult_513_C415_n256), .C(dp_cluster_3_mult_513_C415_n284), 
        .CIX(dp_cluster_3_mult_513_C415_n109), .D(
        dp_cluster_3_mult_513_C415_n312), .CO(dp_cluster_3_mult_513_C415_n104), 
        .COX(dp_cluster_3_mult_513_C415_n103), .S(
        dp_cluster_3_mult_513_C415_n105) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U89 ( .A(dp_cluster_3_mult_513_C415_n112), .B(dp_cluster_3_mult_513_C415_n270), .C(dp_cluster_3_mult_513_C415_n105), 
        .CIX(dp_cluster_3_mult_513_C415_n106), .D(
        dp_cluster_3_mult_513_C415_n110), .CO(dp_cluster_3_mult_513_C415_n101), 
        .COX(dp_cluster_3_mult_513_C415_n100), .S(
        dp_cluster_3_mult_513_C415_n102) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U86 ( .A(dp_cluster_3_mult_513_C415_n103), .B(dp_cluster_3_mult_513_C415_n283), .C(dp_cluster_3_mult_513_C415_n97), 
        .CIX(dp_cluster_3_mult_513_C415_n100), .D(
        dp_cluster_3_mult_513_C415_n104), .CO(dp_cluster_3_mult_513_C415_n94), 
        .COX(dp_cluster_3_mult_513_C415_n93), .S(
        dp_cluster_3_mult_513_C415_n95) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U84 ( .A(dp_cluster_3_mult_513_C415_n98), 
        .B(dp_cluster_3_mult_513_C415_n282), .C(dp_cluster_3_mult_513_C415_n96), .CIX(dp_cluster_3_mult_513_C415_n93), .D(dp_cluster_3_mult_513_C415_n92), 
        .CO(dp_cluster_3_mult_513_C415_n89), .COX(
        dp_cluster_3_mult_513_C415_n88), .S(dp_cluster_3_mult_513_C415_n90) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U82 ( .A(dp_cluster_3_mult_513_C415_n253), .B(dp_cluster_3_mult_513_C415_n267), .C(n1260), .CIX(
        dp_cluster_3_mult_513_C415_n88), .D(dp_cluster_3_mult_513_C415_n91), 
        .CO(dp_cluster_3_mult_513_C415_n84), .COX(
        dp_cluster_3_mult_513_C415_n83), .S(dp_cluster_3_mult_513_C415_n85) );
  CMPE42D1 dp_cluster_3_mult_513_C415_U81 ( .A(dp_cluster_3_mult_513_C415_n266), .B(dp_cluster_3_mult_513_C415_n86), .C(dp_cluster_3_mult_513_C415_n252), 
        .CIX(dp_cluster_3_mult_513_C415_n83), .D(
        dp_cluster_3_mult_513_C415_n281), .CO(dp_cluster_3_mult_513_C415_n81), 
        .COX(dp_cluster_3_mult_513_C415_n80), .S(
        dp_cluster_3_mult_513_C415_n82) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U139 ( .A(
        dp_cluster_2_mult_485_C409_n371), .B(dp_cluster_2_mult_485_C409_n328), 
        .C(dp_cluster_2_mult_485_C409_n342), .CIX(
        dp_cluster_2_mult_485_C409_n237), .D(dp_cluster_2_mult_485_C409_n356), 
        .CO(dp_cluster_2_mult_485_C409_n233), .COX(
        dp_cluster_2_mult_485_C409_n232), .S(dp_cluster_2_mult_485_C409_n234)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U137 ( .A(
        dp_cluster_2_mult_485_C409_n341), .B(dp_cluster_2_mult_485_C409_n370), 
        .C(dp_cluster_2_mult_485_C409_n355), .CIX(
        dp_cluster_2_mult_485_C409_n232), .D(dp_cluster_2_mult_485_C409_n231), 
        .CO(dp_cluster_2_mult_485_C409_n228), .COX(
        dp_cluster_2_mult_485_C409_n227), .S(dp_cluster_2_mult_485_C409_n229)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U135 ( .A(
        dp_cluster_2_mult_485_C409_n354), .B(dp_cluster_2_mult_485_C409_n369), 
        .C(dp_cluster_2_mult_485_C409_n230), .CIX(
        dp_cluster_2_mult_485_C409_n226), .D(dp_cluster_2_mult_485_C409_n227), 
        .CO(dp_cluster_2_mult_485_C409_n223), .COX(
        dp_cluster_2_mult_485_C409_n222), .S(dp_cluster_2_mult_485_C409_n224)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U132 ( .A(
        dp_cluster_2_mult_485_C409_n221), .B(dp_cluster_2_mult_485_C409_n368), 
        .C(dp_cluster_2_mult_485_C409_n225), .CIX(
        dp_cluster_2_mult_485_C409_n222), .D(dp_cluster_2_mult_485_C409_n219), 
        .CO(dp_cluster_2_mult_485_C409_n216), .COX(
        dp_cluster_2_mult_485_C409_n215), .S(dp_cluster_2_mult_485_C409_n217)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U131 ( .A(
        dp_cluster_2_mult_485_C409_n324), .B(dp_cluster_2_mult_485_C409_n295), 
        .C(dp_cluster_2_mult_485_C409_n309), .CIX(
        dp_cluster_2_mult_485_C409_n220), .D(dp_cluster_2_mult_485_C409_n338), 
        .CO(dp_cluster_2_mult_485_C409_n213), .COX(
        dp_cluster_2_mult_485_C409_n212), .S(dp_cluster_2_mult_485_C409_n214)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U130 ( .A(
        dp_cluster_2_mult_485_C409_n352), .B(dp_cluster_2_mult_485_C409_n367), 
        .C(dp_cluster_2_mult_485_C409_n218), .CIX(
        dp_cluster_2_mult_485_C409_n214), .D(dp_cluster_2_mult_485_C409_n215), 
        .CO(dp_cluster_2_mult_485_C409_n210), .COX(
        dp_cluster_2_mult_485_C409_n209), .S(dp_cluster_2_mult_485_C409_n211)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U128 ( .A(
        dp_cluster_2_mult_485_C409_n366), .B(dp_cluster_2_mult_485_C409_n337), 
        .C(dp_cluster_2_mult_485_C409_n351), .CIX(
        dp_cluster_2_mult_485_C409_n212), .D(dp_cluster_2_mult_485_C409_n308), 
        .CO(dp_cluster_2_mult_485_C409_n205), .COX(
        dp_cluster_2_mult_485_C409_n204), .S(dp_cluster_2_mult_485_C409_n206)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U127 ( .A(
        dp_cluster_2_mult_485_C409_n208), .B(dp_cluster_2_mult_485_C409_n323), 
        .C(dp_cluster_2_mult_485_C409_n209), .CIX(
        dp_cluster_2_mult_485_C409_n213), .D(dp_cluster_2_mult_485_C409_n206), 
        .CO(dp_cluster_2_mult_485_C409_n202), .COX(
        dp_cluster_2_mult_485_C409_n201), .S(dp_cluster_2_mult_485_C409_n203)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U125 ( .A(
        dp_cluster_2_mult_485_C409_n322), .B(dp_cluster_2_mult_485_C409_n365), 
        .C(dp_cluster_2_mult_485_C409_n350), .CIX(
        dp_cluster_2_mult_485_C409_n200), .D(dp_cluster_2_mult_485_C409_n207), 
        .CO(dp_cluster_2_mult_485_C409_n197), .COX(
        dp_cluster_2_mult_485_C409_n196), .S(dp_cluster_2_mult_485_C409_n198)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U124 ( .A(
        dp_cluster_2_mult_485_C409_n204), .B(dp_cluster_2_mult_485_C409_n336), 
        .C(dp_cluster_2_mult_485_C409_n198), .CIX(
        dp_cluster_2_mult_485_C409_n201), .D(dp_cluster_2_mult_485_C409_n205), 
        .CO(dp_cluster_2_mult_485_C409_n194), .COX(
        dp_cluster_2_mult_485_C409_n193), .S(dp_cluster_2_mult_485_C409_n195)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U121 ( .A(
        dp_cluster_2_mult_485_C409_n306), .B(dp_cluster_2_mult_485_C409_n349), 
        .C(dp_cluster_2_mult_485_C409_n335), .CIX(
        dp_cluster_2_mult_485_C409_n190), .D(dp_cluster_2_mult_485_C409_n192), 
        .CO(dp_cluster_2_mult_485_C409_n187), .COX(
        dp_cluster_2_mult_485_C409_n186), .S(dp_cluster_2_mult_485_C409_n188)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U120 ( .A(
        dp_cluster_2_mult_485_C409_n199), .B(dp_cluster_2_mult_485_C409_n196), 
        .C(dp_cluster_2_mult_485_C409_n188), .CIX(
        dp_cluster_2_mult_485_C409_n193), .D(dp_cluster_2_mult_485_C409_n197), 
        .CO(dp_cluster_2_mult_485_C409_n184), .COX(
        dp_cluster_2_mult_485_C409_n183), .S(dp_cluster_2_mult_485_C409_n185)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U119 ( .A(
        dp_cluster_2_mult_485_C409_n291), .B(dp_cluster_2_mult_485_C409_n264), 
        .C(dp_cluster_2_mult_485_C409_n278), .CIX(
        dp_cluster_2_mult_485_C409_n191), .D(dp_cluster_2_mult_485_C409_n305), 
        .CO(dp_cluster_2_mult_485_C409_n181), .COX(
        dp_cluster_2_mult_485_C409_n180), .S(dp_cluster_2_mult_485_C409_n182)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U118 ( .A(
        dp_cluster_2_mult_485_C409_n363), .B(dp_cluster_2_mult_485_C409_n334), 
        .C(dp_cluster_2_mult_485_C409_n348), .CIX(
        dp_cluster_2_mult_485_C409_n189), .D(dp_cluster_2_mult_485_C409_n320), 
        .CO(dp_cluster_2_mult_485_C409_n178), .COX(
        dp_cluster_2_mult_485_C409_n177), .S(dp_cluster_2_mult_485_C409_n179)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U117 ( .A(
        dp_cluster_2_mult_485_C409_n182), .B(dp_cluster_2_mult_485_C409_n186), 
        .C(dp_cluster_2_mult_485_C409_n179), .CIX(
        dp_cluster_2_mult_485_C409_n183), .D(dp_cluster_2_mult_485_C409_n187), 
        .CO(dp_cluster_2_mult_485_C409_n175), .COX(
        dp_cluster_2_mult_485_C409_n174), .S(dp_cluster_2_mult_485_C409_n176)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U115 ( .A(
        dp_cluster_2_mult_485_C409_n362), .B(dp_cluster_2_mult_485_C409_n304), 
        .C(dp_cluster_2_mult_485_C409_n347), .CIX(
        dp_cluster_2_mult_485_C409_n180), .D(dp_cluster_2_mult_485_C409_n333), 
        .CO(dp_cluster_2_mult_485_C409_n170), .COX(
        dp_cluster_2_mult_485_C409_n169), .S(dp_cluster_2_mult_485_C409_n171)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U114 ( .A(
        dp_cluster_2_mult_485_C409_n277), .B(dp_cluster_2_mult_485_C409_n319), 
        .C(dp_cluster_2_mult_485_C409_n290), .CIX(
        dp_cluster_2_mult_485_C409_n177), .D(dp_cluster_2_mult_485_C409_n173), 
        .CO(dp_cluster_2_mult_485_C409_n167), .COX(
        dp_cluster_2_mult_485_C409_n166), .S(dp_cluster_2_mult_485_C409_n168)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U113 ( .A(
        dp_cluster_2_mult_485_C409_n168), .B(dp_cluster_2_mult_485_C409_n171), 
        .C(dp_cluster_2_mult_485_C409_n178), .CIX(
        dp_cluster_2_mult_485_C409_n174), .D(dp_cluster_2_mult_485_C409_n181), 
        .CO(dp_cluster_2_mult_485_C409_n164), .COX(
        dp_cluster_2_mult_485_C409_n163), .S(dp_cluster_2_mult_485_C409_n165)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U110 ( .A(
        dp_cluster_2_mult_485_C409_n262), .B(dp_cluster_2_mult_485_C409_n289), 
        .C(dp_cluster_2_mult_485_C409_n361), .CIX(
        dp_cluster_2_mult_485_C409_n169), .D(dp_cluster_2_mult_485_C409_n172), 
        .CO(dp_cluster_2_mult_485_C409_n159), .COX(
        dp_cluster_2_mult_485_C409_n158), .S(dp_cluster_2_mult_485_C409_n160)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U109 ( .A(
        dp_cluster_2_mult_485_C409_n303), .B(dp_cluster_2_mult_485_C409_n346), 
        .C(dp_cluster_2_mult_485_C409_n332), .CIX(
        dp_cluster_2_mult_485_C409_n166), .D(dp_cluster_2_mult_485_C409_n162), 
        .CO(dp_cluster_2_mult_485_C409_n156), .COX(
        dp_cluster_2_mult_485_C409_n155), .S(dp_cluster_2_mult_485_C409_n157)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U108 ( .A(
        dp_cluster_2_mult_485_C409_n170), .B(dp_cluster_2_mult_485_C409_n160), 
        .C(dp_cluster_2_mult_485_C409_n167), .CIX(
        dp_cluster_2_mult_485_C409_n163), .D(dp_cluster_2_mult_485_C409_n157), 
        .CO(dp_cluster_2_mult_485_C409_n153), .COX(
        dp_cluster_2_mult_485_C409_n152), .S(dp_cluster_2_mult_485_C409_n154)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U106 ( .A(
        dp_cluster_2_mult_485_C409_n331), .B(dp_cluster_2_mult_485_C409_n275), 
        .C(n1131), .CIX(dp_cluster_2_mult_485_C409_n158), .D(
        dp_cluster_2_mult_485_C409_n161), .CO(dp_cluster_2_mult_485_C409_n148), 
        .COX(dp_cluster_2_mult_485_C409_n147), .S(
        dp_cluster_2_mult_485_C409_n149) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U105 ( .A(
        dp_cluster_2_mult_485_C409_n317), .B(dp_cluster_2_mult_485_C409_n288), 
        .C(dp_cluster_2_mult_485_C409_n302), .CIX(
        dp_cluster_2_mult_485_C409_n155), .D(dp_cluster_2_mult_485_C409_n261), 
        .CO(dp_cluster_2_mult_485_C409_n145), .COX(
        dp_cluster_2_mult_485_C409_n144), .S(dp_cluster_2_mult_485_C409_n146)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U104 ( .A(
        dp_cluster_2_mult_485_C409_n149), .B(dp_cluster_2_mult_485_C409_n146), 
        .C(dp_cluster_2_mult_485_C409_n156), .CIX(
        dp_cluster_2_mult_485_C409_n152), .D(dp_cluster_2_mult_485_C409_n159), 
        .CO(dp_cluster_2_mult_485_C409_n142), .COX(
        dp_cluster_2_mult_485_C409_n141), .S(dp_cluster_2_mult_485_C409_n143)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U103 ( .A(
        dp_cluster_2_mult_485_C409_n150), .B(dp_cluster_2_mult_485_C409_n260), 
        .C(dp_cluster_2_mult_485_C409_n274), .CIX(
        dp_cluster_2_mult_485_C409_n147), .D(dp_cluster_2_mult_485_C409_n345), 
        .CO(dp_cluster_2_mult_485_C409_n139), .COX(
        dp_cluster_2_mult_485_C409_n138), .S(dp_cluster_2_mult_485_C409_n140)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U102 ( .A(
        dp_cluster_2_mult_485_C409_n330), .B(dp_cluster_2_mult_485_C409_n301), 
        .C(dp_cluster_2_mult_485_C409_n316), .CIX(
        dp_cluster_2_mult_485_C409_n144), .D(dp_cluster_2_mult_485_C409_n287), 
        .CO(dp_cluster_2_mult_485_C409_n136), .COX(
        dp_cluster_2_mult_485_C409_n135), .S(dp_cluster_2_mult_485_C409_n137)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U101 ( .A(
        dp_cluster_2_mult_485_C409_n140), .B(dp_cluster_2_mult_485_C409_n137), 
        .C(dp_cluster_2_mult_485_C409_n145), .CIX(
        dp_cluster_2_mult_485_C409_n141), .D(dp_cluster_2_mult_485_C409_n148), 
        .CO(dp_cluster_2_mult_485_C409_n133), .COX(
        dp_cluster_2_mult_485_C409_n132), .S(dp_cluster_2_mult_485_C409_n134)
         );
  CMPE42D1 dp_cluster_2_mult_485_C409_U98 ( .A(dp_cluster_2_mult_485_C409_n259), .B(dp_cluster_2_mult_485_C409_n300), .C(dp_cluster_2_mult_485_C409_n286), 
        .CIX(dp_cluster_2_mult_485_C409_n129), .D(
        dp_cluster_2_mult_485_C409_n135), .CO(dp_cluster_2_mult_485_C409_n126), 
        .COX(dp_cluster_2_mult_485_C409_n125), .S(
        dp_cluster_2_mult_485_C409_n127) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U97 ( .A(dp_cluster_2_mult_485_C409_n139), .B(dp_cluster_2_mult_485_C409_n138), .C(dp_cluster_2_mult_485_C409_n136), 
        .CIX(dp_cluster_2_mult_485_C409_n132), .D(
        dp_cluster_2_mult_485_C409_n127), .CO(dp_cluster_2_mult_485_C409_n123), 
        .COX(dp_cluster_2_mult_485_C409_n122), .S(
        dp_cluster_2_mult_485_C409_n124) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U95 ( .A(dp_cluster_2_mult_485_C409_n314), .B(dp_cluster_2_mult_485_C409_n285), .C(dp_cluster_2_mult_485_C409_n299), 
        .CIX(dp_cluster_2_mult_485_C409_n121), .D(
        dp_cluster_2_mult_485_C409_n272), .CO(dp_cluster_2_mult_485_C409_n118), 
        .COX(dp_cluster_2_mult_485_C409_n117), .S(
        dp_cluster_2_mult_485_C409_n119) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U94 ( .A(dp_cluster_2_mult_485_C409_n128), .B(dp_cluster_2_mult_485_C409_n125), .C(dp_cluster_2_mult_485_C409_n119), 
        .CIX(dp_cluster_2_mult_485_C409_n122), .D(
        dp_cluster_2_mult_485_C409_n126), .CO(dp_cluster_2_mult_485_C409_n115), 
        .COX(dp_cluster_2_mult_485_C409_n114), .S(
        dp_cluster_2_mult_485_C409_n116) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U92 ( .A(dp_cluster_2_mult_485_C409_n313), .B(dp_cluster_2_mult_485_C409_n271), .C(dp_cluster_2_mult_485_C409_n298), 
        .CIX(dp_cluster_2_mult_485_C409_n120), .D(n1115), .CO(
        dp_cluster_2_mult_485_C409_n110), .COX(dp_cluster_2_mult_485_C409_n109), .S(dp_cluster_2_mult_485_C409_n111) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U91 ( .A(dp_cluster_2_mult_485_C409_n117), .B(dp_cluster_2_mult_485_C409_n257), .C(dp_cluster_2_mult_485_C409_n111), 
        .CIX(dp_cluster_2_mult_485_C409_n114), .D(
        dp_cluster_2_mult_485_C409_n118), .CO(dp_cluster_2_mult_485_C409_n107), 
        .COX(dp_cluster_2_mult_485_C409_n106), .S(
        dp_cluster_2_mult_485_C409_n108) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U90 ( .A(dp_cluster_2_mult_485_C409_n297), .B(dp_cluster_2_mult_485_C409_n256), .C(dp_cluster_2_mult_485_C409_n284), 
        .CIX(dp_cluster_2_mult_485_C409_n109), .D(
        dp_cluster_2_mult_485_C409_n312), .CO(dp_cluster_2_mult_485_C409_n104), 
        .COX(dp_cluster_2_mult_485_C409_n103), .S(
        dp_cluster_2_mult_485_C409_n105) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U89 ( .A(dp_cluster_2_mult_485_C409_n112), .B(dp_cluster_2_mult_485_C409_n270), .C(dp_cluster_2_mult_485_C409_n105), 
        .CIX(dp_cluster_2_mult_485_C409_n106), .D(
        dp_cluster_2_mult_485_C409_n110), .CO(dp_cluster_2_mult_485_C409_n101), 
        .COX(dp_cluster_2_mult_485_C409_n100), .S(
        dp_cluster_2_mult_485_C409_n102) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U86 ( .A(dp_cluster_2_mult_485_C409_n103), .B(dp_cluster_2_mult_485_C409_n283), .C(dp_cluster_2_mult_485_C409_n97), 
        .CIX(dp_cluster_2_mult_485_C409_n100), .D(
        dp_cluster_2_mult_485_C409_n104), .CO(dp_cluster_2_mult_485_C409_n94), 
        .COX(dp_cluster_2_mult_485_C409_n93), .S(
        dp_cluster_2_mult_485_C409_n95) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U84 ( .A(dp_cluster_2_mult_485_C409_n98), 
        .B(dp_cluster_2_mult_485_C409_n282), .C(dp_cluster_2_mult_485_C409_n96), .CIX(dp_cluster_2_mult_485_C409_n93), .D(dp_cluster_2_mult_485_C409_n92), 
        .CO(dp_cluster_2_mult_485_C409_n89), .COX(
        dp_cluster_2_mult_485_C409_n88), .S(dp_cluster_2_mult_485_C409_n90) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U82 ( .A(dp_cluster_2_mult_485_C409_n253), .B(dp_cluster_2_mult_485_C409_n267), .C(n1117), .CIX(
        dp_cluster_2_mult_485_C409_n88), .D(dp_cluster_2_mult_485_C409_n91), 
        .CO(dp_cluster_2_mult_485_C409_n84), .COX(
        dp_cluster_2_mult_485_C409_n83), .S(dp_cluster_2_mult_485_C409_n85) );
  CMPE42D1 dp_cluster_2_mult_485_C409_U81 ( .A(dp_cluster_2_mult_485_C409_n266), .B(dp_cluster_2_mult_485_C409_n86), .C(dp_cluster_2_mult_485_C409_n252), 
        .CIX(dp_cluster_2_mult_485_C409_n83), .D(
        dp_cluster_2_mult_485_C409_n281), .CO(dp_cluster_2_mult_485_C409_n81), 
        .COX(dp_cluster_2_mult_485_C409_n80), .S(
        dp_cluster_2_mult_485_C409_n82) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U139 ( .A(
        dp_cluster_2_mult_486_C409_n371), .B(dp_cluster_2_mult_486_C409_n328), 
        .C(dp_cluster_2_mult_486_C409_n342), .CIX(
        dp_cluster_2_mult_486_C409_n237), .D(dp_cluster_2_mult_486_C409_n356), 
        .CO(dp_cluster_2_mult_486_C409_n233), .COX(
        dp_cluster_2_mult_486_C409_n232), .S(dp_cluster_2_mult_486_C409_n234)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U137 ( .A(
        dp_cluster_2_mult_486_C409_n341), .B(dp_cluster_2_mult_486_C409_n370), 
        .C(dp_cluster_2_mult_486_C409_n355), .CIX(
        dp_cluster_2_mult_486_C409_n232), .D(dp_cluster_2_mult_486_C409_n231), 
        .CO(dp_cluster_2_mult_486_C409_n228), .COX(
        dp_cluster_2_mult_486_C409_n227), .S(dp_cluster_2_mult_486_C409_n229)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U135 ( .A(
        dp_cluster_2_mult_486_C409_n354), .B(dp_cluster_2_mult_486_C409_n369), 
        .C(dp_cluster_2_mult_486_C409_n230), .CIX(
        dp_cluster_2_mult_486_C409_n226), .D(dp_cluster_2_mult_486_C409_n227), 
        .CO(dp_cluster_2_mult_486_C409_n223), .COX(
        dp_cluster_2_mult_486_C409_n222), .S(dp_cluster_2_mult_486_C409_n224)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U132 ( .A(
        dp_cluster_2_mult_486_C409_n221), .B(dp_cluster_2_mult_486_C409_n368), 
        .C(dp_cluster_2_mult_486_C409_n225), .CIX(
        dp_cluster_2_mult_486_C409_n222), .D(dp_cluster_2_mult_486_C409_n219), 
        .CO(dp_cluster_2_mult_486_C409_n216), .COX(
        dp_cluster_2_mult_486_C409_n215), .S(dp_cluster_2_mult_486_C409_n217)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U131 ( .A(
        dp_cluster_2_mult_486_C409_n324), .B(dp_cluster_2_mult_486_C409_n295), 
        .C(dp_cluster_2_mult_486_C409_n309), .CIX(
        dp_cluster_2_mult_486_C409_n220), .D(dp_cluster_2_mult_486_C409_n338), 
        .CO(dp_cluster_2_mult_486_C409_n213), .COX(
        dp_cluster_2_mult_486_C409_n212), .S(dp_cluster_2_mult_486_C409_n214)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U130 ( .A(
        dp_cluster_2_mult_486_C409_n352), .B(dp_cluster_2_mult_486_C409_n367), 
        .C(dp_cluster_2_mult_486_C409_n218), .CIX(
        dp_cluster_2_mult_486_C409_n214), .D(dp_cluster_2_mult_486_C409_n215), 
        .CO(dp_cluster_2_mult_486_C409_n210), .COX(
        dp_cluster_2_mult_486_C409_n209), .S(dp_cluster_2_mult_486_C409_n211)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U128 ( .A(
        dp_cluster_2_mult_486_C409_n366), .B(dp_cluster_2_mult_486_C409_n337), 
        .C(dp_cluster_2_mult_486_C409_n351), .CIX(
        dp_cluster_2_mult_486_C409_n212), .D(dp_cluster_2_mult_486_C409_n308), 
        .CO(dp_cluster_2_mult_486_C409_n205), .COX(
        dp_cluster_2_mult_486_C409_n204), .S(dp_cluster_2_mult_486_C409_n206)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U127 ( .A(
        dp_cluster_2_mult_486_C409_n208), .B(dp_cluster_2_mult_486_C409_n323), 
        .C(dp_cluster_2_mult_486_C409_n209), .CIX(
        dp_cluster_2_mult_486_C409_n213), .D(dp_cluster_2_mult_486_C409_n206), 
        .CO(dp_cluster_2_mult_486_C409_n202), .COX(
        dp_cluster_2_mult_486_C409_n201), .S(dp_cluster_2_mult_486_C409_n203)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U125 ( .A(
        dp_cluster_2_mult_486_C409_n322), .B(dp_cluster_2_mult_486_C409_n365), 
        .C(dp_cluster_2_mult_486_C409_n350), .CIX(
        dp_cluster_2_mult_486_C409_n200), .D(dp_cluster_2_mult_486_C409_n207), 
        .CO(dp_cluster_2_mult_486_C409_n197), .COX(
        dp_cluster_2_mult_486_C409_n196), .S(dp_cluster_2_mult_486_C409_n198)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U124 ( .A(
        dp_cluster_2_mult_486_C409_n204), .B(dp_cluster_2_mult_486_C409_n336), 
        .C(dp_cluster_2_mult_486_C409_n198), .CIX(
        dp_cluster_2_mult_486_C409_n201), .D(dp_cluster_2_mult_486_C409_n205), 
        .CO(dp_cluster_2_mult_486_C409_n194), .COX(
        dp_cluster_2_mult_486_C409_n193), .S(dp_cluster_2_mult_486_C409_n195)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U121 ( .A(
        dp_cluster_2_mult_486_C409_n306), .B(dp_cluster_2_mult_486_C409_n349), 
        .C(dp_cluster_2_mult_486_C409_n335), .CIX(
        dp_cluster_2_mult_486_C409_n190), .D(dp_cluster_2_mult_486_C409_n192), 
        .CO(dp_cluster_2_mult_486_C409_n187), .COX(
        dp_cluster_2_mult_486_C409_n186), .S(dp_cluster_2_mult_486_C409_n188)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U120 ( .A(
        dp_cluster_2_mult_486_C409_n199), .B(dp_cluster_2_mult_486_C409_n196), 
        .C(dp_cluster_2_mult_486_C409_n188), .CIX(
        dp_cluster_2_mult_486_C409_n193), .D(dp_cluster_2_mult_486_C409_n197), 
        .CO(dp_cluster_2_mult_486_C409_n184), .COX(
        dp_cluster_2_mult_486_C409_n183), .S(dp_cluster_2_mult_486_C409_n185)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U119 ( .A(
        dp_cluster_2_mult_486_C409_n291), .B(dp_cluster_2_mult_486_C409_n264), 
        .C(dp_cluster_2_mult_486_C409_n278), .CIX(
        dp_cluster_2_mult_486_C409_n191), .D(dp_cluster_2_mult_486_C409_n305), 
        .CO(dp_cluster_2_mult_486_C409_n181), .COX(
        dp_cluster_2_mult_486_C409_n180), .S(dp_cluster_2_mult_486_C409_n182)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U118 ( .A(
        dp_cluster_2_mult_486_C409_n363), .B(dp_cluster_2_mult_486_C409_n334), 
        .C(dp_cluster_2_mult_486_C409_n348), .CIX(
        dp_cluster_2_mult_486_C409_n189), .D(dp_cluster_2_mult_486_C409_n320), 
        .CO(dp_cluster_2_mult_486_C409_n178), .COX(
        dp_cluster_2_mult_486_C409_n177), .S(dp_cluster_2_mult_486_C409_n179)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U117 ( .A(
        dp_cluster_2_mult_486_C409_n182), .B(dp_cluster_2_mult_486_C409_n186), 
        .C(dp_cluster_2_mult_486_C409_n179), .CIX(
        dp_cluster_2_mult_486_C409_n183), .D(dp_cluster_2_mult_486_C409_n187), 
        .CO(dp_cluster_2_mult_486_C409_n175), .COX(
        dp_cluster_2_mult_486_C409_n174), .S(dp_cluster_2_mult_486_C409_n176)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U115 ( .A(
        dp_cluster_2_mult_486_C409_n362), .B(dp_cluster_2_mult_486_C409_n304), 
        .C(dp_cluster_2_mult_486_C409_n347), .CIX(
        dp_cluster_2_mult_486_C409_n180), .D(dp_cluster_2_mult_486_C409_n333), 
        .CO(dp_cluster_2_mult_486_C409_n170), .COX(
        dp_cluster_2_mult_486_C409_n169), .S(dp_cluster_2_mult_486_C409_n171)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U114 ( .A(
        dp_cluster_2_mult_486_C409_n277), .B(dp_cluster_2_mult_486_C409_n319), 
        .C(dp_cluster_2_mult_486_C409_n290), .CIX(
        dp_cluster_2_mult_486_C409_n177), .D(dp_cluster_2_mult_486_C409_n173), 
        .CO(dp_cluster_2_mult_486_C409_n167), .COX(
        dp_cluster_2_mult_486_C409_n166), .S(dp_cluster_2_mult_486_C409_n168)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U113 ( .A(
        dp_cluster_2_mult_486_C409_n168), .B(dp_cluster_2_mult_486_C409_n171), 
        .C(dp_cluster_2_mult_486_C409_n178), .CIX(
        dp_cluster_2_mult_486_C409_n174), .D(dp_cluster_2_mult_486_C409_n181), 
        .CO(dp_cluster_2_mult_486_C409_n164), .COX(
        dp_cluster_2_mult_486_C409_n163), .S(dp_cluster_2_mult_486_C409_n165)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U110 ( .A(
        dp_cluster_2_mult_486_C409_n262), .B(dp_cluster_2_mult_486_C409_n289), 
        .C(dp_cluster_2_mult_486_C409_n361), .CIX(
        dp_cluster_2_mult_486_C409_n169), .D(dp_cluster_2_mult_486_C409_n172), 
        .CO(dp_cluster_2_mult_486_C409_n159), .COX(
        dp_cluster_2_mult_486_C409_n158), .S(dp_cluster_2_mult_486_C409_n160)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U109 ( .A(
        dp_cluster_2_mult_486_C409_n303), .B(dp_cluster_2_mult_486_C409_n346), 
        .C(dp_cluster_2_mult_486_C409_n332), .CIX(
        dp_cluster_2_mult_486_C409_n166), .D(dp_cluster_2_mult_486_C409_n162), 
        .CO(dp_cluster_2_mult_486_C409_n156), .COX(
        dp_cluster_2_mult_486_C409_n155), .S(dp_cluster_2_mult_486_C409_n157)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U108 ( .A(
        dp_cluster_2_mult_486_C409_n170), .B(dp_cluster_2_mult_486_C409_n160), 
        .C(dp_cluster_2_mult_486_C409_n167), .CIX(
        dp_cluster_2_mult_486_C409_n163), .D(dp_cluster_2_mult_486_C409_n157), 
        .CO(dp_cluster_2_mult_486_C409_n153), .COX(
        dp_cluster_2_mult_486_C409_n152), .S(dp_cluster_2_mult_486_C409_n154)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U106 ( .A(
        dp_cluster_2_mult_486_C409_n331), .B(dp_cluster_2_mult_486_C409_n275), 
        .C(n1269), .CIX(dp_cluster_2_mult_486_C409_n158), .D(
        dp_cluster_2_mult_486_C409_n161), .CO(dp_cluster_2_mult_486_C409_n148), 
        .COX(dp_cluster_2_mult_486_C409_n147), .S(
        dp_cluster_2_mult_486_C409_n149) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U105 ( .A(
        dp_cluster_2_mult_486_C409_n317), .B(dp_cluster_2_mult_486_C409_n288), 
        .C(dp_cluster_2_mult_486_C409_n302), .CIX(
        dp_cluster_2_mult_486_C409_n155), .D(dp_cluster_2_mult_486_C409_n261), 
        .CO(dp_cluster_2_mult_486_C409_n145), .COX(
        dp_cluster_2_mult_486_C409_n144), .S(dp_cluster_2_mult_486_C409_n146)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U104 ( .A(
        dp_cluster_2_mult_486_C409_n149), .B(dp_cluster_2_mult_486_C409_n146), 
        .C(dp_cluster_2_mult_486_C409_n156), .CIX(
        dp_cluster_2_mult_486_C409_n152), .D(dp_cluster_2_mult_486_C409_n159), 
        .CO(dp_cluster_2_mult_486_C409_n142), .COX(
        dp_cluster_2_mult_486_C409_n141), .S(dp_cluster_2_mult_486_C409_n143)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U103 ( .A(
        dp_cluster_2_mult_486_C409_n150), .B(dp_cluster_2_mult_486_C409_n260), 
        .C(dp_cluster_2_mult_486_C409_n274), .CIX(
        dp_cluster_2_mult_486_C409_n147), .D(dp_cluster_2_mult_486_C409_n345), 
        .CO(dp_cluster_2_mult_486_C409_n139), .COX(
        dp_cluster_2_mult_486_C409_n138), .S(dp_cluster_2_mult_486_C409_n140)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U102 ( .A(
        dp_cluster_2_mult_486_C409_n330), .B(dp_cluster_2_mult_486_C409_n301), 
        .C(dp_cluster_2_mult_486_C409_n316), .CIX(
        dp_cluster_2_mult_486_C409_n144), .D(dp_cluster_2_mult_486_C409_n287), 
        .CO(dp_cluster_2_mult_486_C409_n136), .COX(
        dp_cluster_2_mult_486_C409_n135), .S(dp_cluster_2_mult_486_C409_n137)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U101 ( .A(
        dp_cluster_2_mult_486_C409_n140), .B(dp_cluster_2_mult_486_C409_n137), 
        .C(dp_cluster_2_mult_486_C409_n145), .CIX(
        dp_cluster_2_mult_486_C409_n141), .D(dp_cluster_2_mult_486_C409_n148), 
        .CO(dp_cluster_2_mult_486_C409_n133), .COX(
        dp_cluster_2_mult_486_C409_n132), .S(dp_cluster_2_mult_486_C409_n134)
         );
  CMPE42D1 dp_cluster_2_mult_486_C409_U98 ( .A(dp_cluster_2_mult_486_C409_n259), .B(dp_cluster_2_mult_486_C409_n300), .C(dp_cluster_2_mult_486_C409_n286), 
        .CIX(dp_cluster_2_mult_486_C409_n129), .D(
        dp_cluster_2_mult_486_C409_n135), .CO(dp_cluster_2_mult_486_C409_n126), 
        .COX(dp_cluster_2_mult_486_C409_n125), .S(
        dp_cluster_2_mult_486_C409_n127) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U97 ( .A(dp_cluster_2_mult_486_C409_n139), .B(dp_cluster_2_mult_486_C409_n138), .C(dp_cluster_2_mult_486_C409_n136), 
        .CIX(dp_cluster_2_mult_486_C409_n132), .D(
        dp_cluster_2_mult_486_C409_n127), .CO(dp_cluster_2_mult_486_C409_n123), 
        .COX(dp_cluster_2_mult_486_C409_n122), .S(
        dp_cluster_2_mult_486_C409_n124) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U95 ( .A(dp_cluster_2_mult_486_C409_n314), .B(dp_cluster_2_mult_486_C409_n285), .C(dp_cluster_2_mult_486_C409_n299), 
        .CIX(dp_cluster_2_mult_486_C409_n121), .D(
        dp_cluster_2_mult_486_C409_n272), .CO(dp_cluster_2_mult_486_C409_n118), 
        .COX(dp_cluster_2_mult_486_C409_n117), .S(
        dp_cluster_2_mult_486_C409_n119) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U94 ( .A(dp_cluster_2_mult_486_C409_n128), .B(dp_cluster_2_mult_486_C409_n125), .C(dp_cluster_2_mult_486_C409_n119), 
        .CIX(dp_cluster_2_mult_486_C409_n122), .D(
        dp_cluster_2_mult_486_C409_n126), .CO(dp_cluster_2_mult_486_C409_n115), 
        .COX(dp_cluster_2_mult_486_C409_n114), .S(
        dp_cluster_2_mult_486_C409_n116) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U92 ( .A(dp_cluster_2_mult_486_C409_n313), .B(dp_cluster_2_mult_486_C409_n271), .C(dp_cluster_2_mult_486_C409_n298), 
        .CIX(dp_cluster_2_mult_486_C409_n120), .D(n1257), .CO(
        dp_cluster_2_mult_486_C409_n110), .COX(dp_cluster_2_mult_486_C409_n109), .S(dp_cluster_2_mult_486_C409_n111) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U91 ( .A(dp_cluster_2_mult_486_C409_n117), .B(dp_cluster_2_mult_486_C409_n257), .C(dp_cluster_2_mult_486_C409_n111), 
        .CIX(dp_cluster_2_mult_486_C409_n114), .D(
        dp_cluster_2_mult_486_C409_n118), .CO(dp_cluster_2_mult_486_C409_n107), 
        .COX(dp_cluster_2_mult_486_C409_n106), .S(
        dp_cluster_2_mult_486_C409_n108) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U90 ( .A(dp_cluster_2_mult_486_C409_n297), .B(dp_cluster_2_mult_486_C409_n256), .C(dp_cluster_2_mult_486_C409_n284), 
        .CIX(dp_cluster_2_mult_486_C409_n109), .D(
        dp_cluster_2_mult_486_C409_n312), .CO(dp_cluster_2_mult_486_C409_n104), 
        .COX(dp_cluster_2_mult_486_C409_n103), .S(
        dp_cluster_2_mult_486_C409_n105) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U89 ( .A(dp_cluster_2_mult_486_C409_n112), .B(dp_cluster_2_mult_486_C409_n270), .C(dp_cluster_2_mult_486_C409_n105), 
        .CIX(dp_cluster_2_mult_486_C409_n106), .D(
        dp_cluster_2_mult_486_C409_n110), .CO(dp_cluster_2_mult_486_C409_n101), 
        .COX(dp_cluster_2_mult_486_C409_n100), .S(
        dp_cluster_2_mult_486_C409_n102) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U86 ( .A(dp_cluster_2_mult_486_C409_n103), .B(dp_cluster_2_mult_486_C409_n283), .C(dp_cluster_2_mult_486_C409_n97), 
        .CIX(dp_cluster_2_mult_486_C409_n100), .D(
        dp_cluster_2_mult_486_C409_n104), .CO(dp_cluster_2_mult_486_C409_n94), 
        .COX(dp_cluster_2_mult_486_C409_n93), .S(
        dp_cluster_2_mult_486_C409_n95) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U84 ( .A(dp_cluster_2_mult_486_C409_n98), 
        .B(dp_cluster_2_mult_486_C409_n282), .C(dp_cluster_2_mult_486_C409_n96), .CIX(dp_cluster_2_mult_486_C409_n93), .D(dp_cluster_2_mult_486_C409_n92), 
        .CO(dp_cluster_2_mult_486_C409_n89), .COX(
        dp_cluster_2_mult_486_C409_n88), .S(dp_cluster_2_mult_486_C409_n90) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U82 ( .A(dp_cluster_2_mult_486_C409_n253), .B(dp_cluster_2_mult_486_C409_n267), .C(n1258), .CIX(
        dp_cluster_2_mult_486_C409_n88), .D(dp_cluster_2_mult_486_C409_n91), 
        .CO(dp_cluster_2_mult_486_C409_n84), .COX(
        dp_cluster_2_mult_486_C409_n83), .S(dp_cluster_2_mult_486_C409_n85) );
  CMPE42D1 dp_cluster_2_mult_486_C409_U81 ( .A(dp_cluster_2_mult_486_C409_n266), .B(dp_cluster_2_mult_486_C409_n86), .C(dp_cluster_2_mult_486_C409_n252), 
        .CIX(dp_cluster_2_mult_486_C409_n83), .D(
        dp_cluster_2_mult_486_C409_n281), .CO(dp_cluster_2_mult_486_C409_n81), 
        .COX(dp_cluster_2_mult_486_C409_n80), .S(
        dp_cluster_2_mult_486_C409_n82) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U139 ( .A(
        dp_cluster_1_mult_512_C418_n371), .B(dp_cluster_1_mult_512_C418_n328), 
        .C(dp_cluster_1_mult_512_C418_n342), .CIX(
        dp_cluster_1_mult_512_C418_n237), .D(dp_cluster_1_mult_512_C418_n356), 
        .CO(dp_cluster_1_mult_512_C418_n233), .COX(
        dp_cluster_1_mult_512_C418_n232), .S(dp_cluster_1_mult_512_C418_n234)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U137 ( .A(
        dp_cluster_1_mult_512_C418_n341), .B(dp_cluster_1_mult_512_C418_n370), 
        .C(dp_cluster_1_mult_512_C418_n355), .CIX(
        dp_cluster_1_mult_512_C418_n232), .D(dp_cluster_1_mult_512_C418_n231), 
        .CO(dp_cluster_1_mult_512_C418_n228), .COX(
        dp_cluster_1_mult_512_C418_n227), .S(dp_cluster_1_mult_512_C418_n229)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U135 ( .A(
        dp_cluster_1_mult_512_C418_n354), .B(dp_cluster_1_mult_512_C418_n369), 
        .C(dp_cluster_1_mult_512_C418_n230), .CIX(
        dp_cluster_1_mult_512_C418_n226), .D(dp_cluster_1_mult_512_C418_n227), 
        .CO(dp_cluster_1_mult_512_C418_n223), .COX(
        dp_cluster_1_mult_512_C418_n222), .S(dp_cluster_1_mult_512_C418_n224)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U132 ( .A(
        dp_cluster_1_mult_512_C418_n221), .B(dp_cluster_1_mult_512_C418_n368), 
        .C(dp_cluster_1_mult_512_C418_n225), .CIX(
        dp_cluster_1_mult_512_C418_n222), .D(dp_cluster_1_mult_512_C418_n219), 
        .CO(dp_cluster_1_mult_512_C418_n216), .COX(
        dp_cluster_1_mult_512_C418_n215), .S(dp_cluster_1_mult_512_C418_n217)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U131 ( .A(
        dp_cluster_1_mult_512_C418_n324), .B(dp_cluster_1_mult_512_C418_n295), 
        .C(dp_cluster_1_mult_512_C418_n309), .CIX(
        dp_cluster_1_mult_512_C418_n220), .D(dp_cluster_1_mult_512_C418_n338), 
        .CO(dp_cluster_1_mult_512_C418_n213), .COX(
        dp_cluster_1_mult_512_C418_n212), .S(dp_cluster_1_mult_512_C418_n214)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U130 ( .A(
        dp_cluster_1_mult_512_C418_n352), .B(dp_cluster_1_mult_512_C418_n367), 
        .C(dp_cluster_1_mult_512_C418_n218), .CIX(
        dp_cluster_1_mult_512_C418_n214), .D(dp_cluster_1_mult_512_C418_n215), 
        .CO(dp_cluster_1_mult_512_C418_n210), .COX(
        dp_cluster_1_mult_512_C418_n209), .S(dp_cluster_1_mult_512_C418_n211)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U128 ( .A(
        dp_cluster_1_mult_512_C418_n366), .B(dp_cluster_1_mult_512_C418_n337), 
        .C(dp_cluster_1_mult_512_C418_n351), .CIX(
        dp_cluster_1_mult_512_C418_n212), .D(dp_cluster_1_mult_512_C418_n308), 
        .CO(dp_cluster_1_mult_512_C418_n205), .COX(
        dp_cluster_1_mult_512_C418_n204), .S(dp_cluster_1_mult_512_C418_n206)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U127 ( .A(
        dp_cluster_1_mult_512_C418_n208), .B(dp_cluster_1_mult_512_C418_n323), 
        .C(dp_cluster_1_mult_512_C418_n209), .CIX(
        dp_cluster_1_mult_512_C418_n213), .D(dp_cluster_1_mult_512_C418_n206), 
        .CO(dp_cluster_1_mult_512_C418_n202), .COX(
        dp_cluster_1_mult_512_C418_n201), .S(dp_cluster_1_mult_512_C418_n203)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U125 ( .A(
        dp_cluster_1_mult_512_C418_n322), .B(dp_cluster_1_mult_512_C418_n365), 
        .C(dp_cluster_1_mult_512_C418_n350), .CIX(
        dp_cluster_1_mult_512_C418_n200), .D(dp_cluster_1_mult_512_C418_n207), 
        .CO(dp_cluster_1_mult_512_C418_n197), .COX(
        dp_cluster_1_mult_512_C418_n196), .S(dp_cluster_1_mult_512_C418_n198)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U124 ( .A(
        dp_cluster_1_mult_512_C418_n204), .B(dp_cluster_1_mult_512_C418_n336), 
        .C(dp_cluster_1_mult_512_C418_n198), .CIX(
        dp_cluster_1_mult_512_C418_n201), .D(dp_cluster_1_mult_512_C418_n205), 
        .CO(dp_cluster_1_mult_512_C418_n194), .COX(
        dp_cluster_1_mult_512_C418_n193), .S(dp_cluster_1_mult_512_C418_n195)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U121 ( .A(
        dp_cluster_1_mult_512_C418_n306), .B(dp_cluster_1_mult_512_C418_n349), 
        .C(dp_cluster_1_mult_512_C418_n335), .CIX(
        dp_cluster_1_mult_512_C418_n190), .D(dp_cluster_1_mult_512_C418_n192), 
        .CO(dp_cluster_1_mult_512_C418_n187), .COX(
        dp_cluster_1_mult_512_C418_n186), .S(dp_cluster_1_mult_512_C418_n188)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U120 ( .A(
        dp_cluster_1_mult_512_C418_n199), .B(dp_cluster_1_mult_512_C418_n196), 
        .C(dp_cluster_1_mult_512_C418_n188), .CIX(
        dp_cluster_1_mult_512_C418_n193), .D(dp_cluster_1_mult_512_C418_n197), 
        .CO(dp_cluster_1_mult_512_C418_n184), .COX(
        dp_cluster_1_mult_512_C418_n183), .S(dp_cluster_1_mult_512_C418_n185)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U119 ( .A(
        dp_cluster_1_mult_512_C418_n291), .B(dp_cluster_1_mult_512_C418_n264), 
        .C(dp_cluster_1_mult_512_C418_n278), .CIX(
        dp_cluster_1_mult_512_C418_n191), .D(dp_cluster_1_mult_512_C418_n305), 
        .CO(dp_cluster_1_mult_512_C418_n181), .COX(
        dp_cluster_1_mult_512_C418_n180), .S(dp_cluster_1_mult_512_C418_n182)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U118 ( .A(
        dp_cluster_1_mult_512_C418_n363), .B(dp_cluster_1_mult_512_C418_n334), 
        .C(dp_cluster_1_mult_512_C418_n348), .CIX(
        dp_cluster_1_mult_512_C418_n189), .D(dp_cluster_1_mult_512_C418_n320), 
        .CO(dp_cluster_1_mult_512_C418_n178), .COX(
        dp_cluster_1_mult_512_C418_n177), .S(dp_cluster_1_mult_512_C418_n179)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U117 ( .A(
        dp_cluster_1_mult_512_C418_n182), .B(dp_cluster_1_mult_512_C418_n186), 
        .C(dp_cluster_1_mult_512_C418_n179), .CIX(
        dp_cluster_1_mult_512_C418_n183), .D(dp_cluster_1_mult_512_C418_n187), 
        .CO(dp_cluster_1_mult_512_C418_n175), .COX(
        dp_cluster_1_mult_512_C418_n174), .S(dp_cluster_1_mult_512_C418_n176)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U115 ( .A(
        dp_cluster_1_mult_512_C418_n362), .B(dp_cluster_1_mult_512_C418_n304), 
        .C(dp_cluster_1_mult_512_C418_n347), .CIX(
        dp_cluster_1_mult_512_C418_n180), .D(dp_cluster_1_mult_512_C418_n333), 
        .CO(dp_cluster_1_mult_512_C418_n170), .COX(
        dp_cluster_1_mult_512_C418_n169), .S(dp_cluster_1_mult_512_C418_n171)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U114 ( .A(
        dp_cluster_1_mult_512_C418_n277), .B(dp_cluster_1_mult_512_C418_n319), 
        .C(dp_cluster_1_mult_512_C418_n290), .CIX(
        dp_cluster_1_mult_512_C418_n177), .D(dp_cluster_1_mult_512_C418_n173), 
        .CO(dp_cluster_1_mult_512_C418_n167), .COX(
        dp_cluster_1_mult_512_C418_n166), .S(dp_cluster_1_mult_512_C418_n168)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U113 ( .A(
        dp_cluster_1_mult_512_C418_n168), .B(dp_cluster_1_mult_512_C418_n171), 
        .C(dp_cluster_1_mult_512_C418_n178), .CIX(
        dp_cluster_1_mult_512_C418_n174), .D(dp_cluster_1_mult_512_C418_n181), 
        .CO(dp_cluster_1_mult_512_C418_n164), .COX(
        dp_cluster_1_mult_512_C418_n163), .S(dp_cluster_1_mult_512_C418_n165)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U110 ( .A(
        dp_cluster_1_mult_512_C418_n262), .B(dp_cluster_1_mult_512_C418_n289), 
        .C(dp_cluster_1_mult_512_C418_n361), .CIX(
        dp_cluster_1_mult_512_C418_n169), .D(dp_cluster_1_mult_512_C418_n172), 
        .CO(dp_cluster_1_mult_512_C418_n159), .COX(
        dp_cluster_1_mult_512_C418_n158), .S(dp_cluster_1_mult_512_C418_n160)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U109 ( .A(
        dp_cluster_1_mult_512_C418_n303), .B(dp_cluster_1_mult_512_C418_n346), 
        .C(dp_cluster_1_mult_512_C418_n332), .CIX(
        dp_cluster_1_mult_512_C418_n166), .D(dp_cluster_1_mult_512_C418_n162), 
        .CO(dp_cluster_1_mult_512_C418_n156), .COX(
        dp_cluster_1_mult_512_C418_n155), .S(dp_cluster_1_mult_512_C418_n157)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U108 ( .A(
        dp_cluster_1_mult_512_C418_n170), .B(dp_cluster_1_mult_512_C418_n160), 
        .C(dp_cluster_1_mult_512_C418_n167), .CIX(
        dp_cluster_1_mult_512_C418_n163), .D(dp_cluster_1_mult_512_C418_n157), 
        .CO(dp_cluster_1_mult_512_C418_n153), .COX(
        dp_cluster_1_mult_512_C418_n152), .S(dp_cluster_1_mult_512_C418_n154)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U106 ( .A(
        dp_cluster_1_mult_512_C418_n331), .B(dp_cluster_1_mult_512_C418_n275), 
        .C(n1172), .CIX(dp_cluster_1_mult_512_C418_n158), .D(
        dp_cluster_1_mult_512_C418_n161), .CO(dp_cluster_1_mult_512_C418_n148), 
        .COX(dp_cluster_1_mult_512_C418_n147), .S(
        dp_cluster_1_mult_512_C418_n149) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U105 ( .A(
        dp_cluster_1_mult_512_C418_n317), .B(dp_cluster_1_mult_512_C418_n288), 
        .C(dp_cluster_1_mult_512_C418_n302), .CIX(
        dp_cluster_1_mult_512_C418_n155), .D(dp_cluster_1_mult_512_C418_n261), 
        .CO(dp_cluster_1_mult_512_C418_n145), .COX(
        dp_cluster_1_mult_512_C418_n144), .S(dp_cluster_1_mult_512_C418_n146)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U104 ( .A(
        dp_cluster_1_mult_512_C418_n149), .B(dp_cluster_1_mult_512_C418_n146), 
        .C(dp_cluster_1_mult_512_C418_n156), .CIX(
        dp_cluster_1_mult_512_C418_n152), .D(dp_cluster_1_mult_512_C418_n159), 
        .CO(dp_cluster_1_mult_512_C418_n142), .COX(
        dp_cluster_1_mult_512_C418_n141), .S(dp_cluster_1_mult_512_C418_n143)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U103 ( .A(
        dp_cluster_1_mult_512_C418_n150), .B(dp_cluster_1_mult_512_C418_n260), 
        .C(dp_cluster_1_mult_512_C418_n274), .CIX(
        dp_cluster_1_mult_512_C418_n147), .D(dp_cluster_1_mult_512_C418_n345), 
        .CO(dp_cluster_1_mult_512_C418_n139), .COX(
        dp_cluster_1_mult_512_C418_n138), .S(dp_cluster_1_mult_512_C418_n140)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U102 ( .A(
        dp_cluster_1_mult_512_C418_n330), .B(dp_cluster_1_mult_512_C418_n301), 
        .C(dp_cluster_1_mult_512_C418_n316), .CIX(
        dp_cluster_1_mult_512_C418_n144), .D(dp_cluster_1_mult_512_C418_n287), 
        .CO(dp_cluster_1_mult_512_C418_n136), .COX(
        dp_cluster_1_mult_512_C418_n135), .S(dp_cluster_1_mult_512_C418_n137)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U101 ( .A(
        dp_cluster_1_mult_512_C418_n140), .B(dp_cluster_1_mult_512_C418_n137), 
        .C(dp_cluster_1_mult_512_C418_n145), .CIX(
        dp_cluster_1_mult_512_C418_n141), .D(dp_cluster_1_mult_512_C418_n148), 
        .CO(dp_cluster_1_mult_512_C418_n133), .COX(
        dp_cluster_1_mult_512_C418_n132), .S(dp_cluster_1_mult_512_C418_n134)
         );
  CMPE42D1 dp_cluster_1_mult_512_C418_U98 ( .A(dp_cluster_1_mult_512_C418_n259), .B(dp_cluster_1_mult_512_C418_n300), .C(dp_cluster_1_mult_512_C418_n286), 
        .CIX(dp_cluster_1_mult_512_C418_n129), .D(
        dp_cluster_1_mult_512_C418_n135), .CO(dp_cluster_1_mult_512_C418_n126), 
        .COX(dp_cluster_1_mult_512_C418_n125), .S(
        dp_cluster_1_mult_512_C418_n127) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U97 ( .A(dp_cluster_1_mult_512_C418_n139), .B(dp_cluster_1_mult_512_C418_n138), .C(dp_cluster_1_mult_512_C418_n136), 
        .CIX(dp_cluster_1_mult_512_C418_n132), .D(
        dp_cluster_1_mult_512_C418_n127), .CO(dp_cluster_1_mult_512_C418_n123), 
        .COX(dp_cluster_1_mult_512_C418_n122), .S(
        dp_cluster_1_mult_512_C418_n124) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U95 ( .A(dp_cluster_1_mult_512_C418_n314), .B(dp_cluster_1_mult_512_C418_n285), .C(dp_cluster_1_mult_512_C418_n299), 
        .CIX(dp_cluster_1_mult_512_C418_n121), .D(
        dp_cluster_1_mult_512_C418_n272), .CO(dp_cluster_1_mult_512_C418_n118), 
        .COX(dp_cluster_1_mult_512_C418_n117), .S(
        dp_cluster_1_mult_512_C418_n119) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U94 ( .A(dp_cluster_1_mult_512_C418_n128), .B(dp_cluster_1_mult_512_C418_n125), .C(dp_cluster_1_mult_512_C418_n119), 
        .CIX(dp_cluster_1_mult_512_C418_n122), .D(
        dp_cluster_1_mult_512_C418_n126), .CO(dp_cluster_1_mult_512_C418_n115), 
        .COX(dp_cluster_1_mult_512_C418_n114), .S(
        dp_cluster_1_mult_512_C418_n116) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U92 ( .A(dp_cluster_1_mult_512_C418_n313), .B(dp_cluster_1_mult_512_C418_n271), .C(dp_cluster_1_mult_512_C418_n298), 
        .CIX(dp_cluster_1_mult_512_C418_n120), .D(n1157), .CO(
        dp_cluster_1_mult_512_C418_n110), .COX(dp_cluster_1_mult_512_C418_n109), .S(dp_cluster_1_mult_512_C418_n111) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U91 ( .A(dp_cluster_1_mult_512_C418_n117), .B(dp_cluster_1_mult_512_C418_n257), .C(dp_cluster_1_mult_512_C418_n111), 
        .CIX(dp_cluster_1_mult_512_C418_n114), .D(
        dp_cluster_1_mult_512_C418_n118), .CO(dp_cluster_1_mult_512_C418_n107), 
        .COX(dp_cluster_1_mult_512_C418_n106), .S(
        dp_cluster_1_mult_512_C418_n108) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U90 ( .A(dp_cluster_1_mult_512_C418_n297), .B(dp_cluster_1_mult_512_C418_n256), .C(dp_cluster_1_mult_512_C418_n284), 
        .CIX(dp_cluster_1_mult_512_C418_n109), .D(
        dp_cluster_1_mult_512_C418_n312), .CO(dp_cluster_1_mult_512_C418_n104), 
        .COX(dp_cluster_1_mult_512_C418_n103), .S(
        dp_cluster_1_mult_512_C418_n105) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U89 ( .A(dp_cluster_1_mult_512_C418_n112), .B(dp_cluster_1_mult_512_C418_n270), .C(dp_cluster_1_mult_512_C418_n105), 
        .CIX(dp_cluster_1_mult_512_C418_n106), .D(
        dp_cluster_1_mult_512_C418_n110), .CO(dp_cluster_1_mult_512_C418_n101), 
        .COX(dp_cluster_1_mult_512_C418_n100), .S(
        dp_cluster_1_mult_512_C418_n102) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U86 ( .A(dp_cluster_1_mult_512_C418_n103), .B(dp_cluster_1_mult_512_C418_n283), .C(dp_cluster_1_mult_512_C418_n97), 
        .CIX(dp_cluster_1_mult_512_C418_n100), .D(
        dp_cluster_1_mult_512_C418_n104), .CO(dp_cluster_1_mult_512_C418_n94), 
        .COX(dp_cluster_1_mult_512_C418_n93), .S(
        dp_cluster_1_mult_512_C418_n95) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U84 ( .A(dp_cluster_1_mult_512_C418_n98), 
        .B(dp_cluster_1_mult_512_C418_n282), .C(dp_cluster_1_mult_512_C418_n96), .CIX(dp_cluster_1_mult_512_C418_n93), .D(dp_cluster_1_mult_512_C418_n92), 
        .CO(dp_cluster_1_mult_512_C418_n89), .COX(
        dp_cluster_1_mult_512_C418_n88), .S(dp_cluster_1_mult_512_C418_n90) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U82 ( .A(dp_cluster_1_mult_512_C418_n253), .B(dp_cluster_1_mult_512_C418_n267), .C(n1158), .CIX(
        dp_cluster_1_mult_512_C418_n88), .D(dp_cluster_1_mult_512_C418_n91), 
        .CO(dp_cluster_1_mult_512_C418_n84), .COX(
        dp_cluster_1_mult_512_C418_n83), .S(dp_cluster_1_mult_512_C418_n85) );
  CMPE42D1 dp_cluster_1_mult_512_C418_U81 ( .A(dp_cluster_1_mult_512_C418_n266), .B(dp_cluster_1_mult_512_C418_n86), .C(dp_cluster_1_mult_512_C418_n252), 
        .CIX(dp_cluster_1_mult_512_C418_n83), .D(
        dp_cluster_1_mult_512_C418_n281), .CO(dp_cluster_1_mult_512_C418_n81), 
        .COX(dp_cluster_1_mult_512_C418_n80), .S(
        dp_cluster_1_mult_512_C418_n82) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U139 ( .A(
        dp_cluster_1_mult_513_C418_n371), .B(dp_cluster_1_mult_513_C418_n328), 
        .C(dp_cluster_1_mult_513_C418_n342), .CIX(
        dp_cluster_1_mult_513_C418_n237), .D(dp_cluster_1_mult_513_C418_n356), 
        .CO(dp_cluster_1_mult_513_C418_n233), .COX(
        dp_cluster_1_mult_513_C418_n232), .S(dp_cluster_1_mult_513_C418_n234)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U137 ( .A(
        dp_cluster_1_mult_513_C418_n341), .B(dp_cluster_1_mult_513_C418_n370), 
        .C(dp_cluster_1_mult_513_C418_n355), .CIX(
        dp_cluster_1_mult_513_C418_n232), .D(dp_cluster_1_mult_513_C418_n231), 
        .CO(dp_cluster_1_mult_513_C418_n228), .COX(
        dp_cluster_1_mult_513_C418_n227), .S(dp_cluster_1_mult_513_C418_n229)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U135 ( .A(
        dp_cluster_1_mult_513_C418_n354), .B(dp_cluster_1_mult_513_C418_n369), 
        .C(dp_cluster_1_mult_513_C418_n230), .CIX(
        dp_cluster_1_mult_513_C418_n226), .D(dp_cluster_1_mult_513_C418_n227), 
        .CO(dp_cluster_1_mult_513_C418_n223), .COX(
        dp_cluster_1_mult_513_C418_n222), .S(dp_cluster_1_mult_513_C418_n224)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U132 ( .A(
        dp_cluster_1_mult_513_C418_n221), .B(dp_cluster_1_mult_513_C418_n368), 
        .C(dp_cluster_1_mult_513_C418_n225), .CIX(
        dp_cluster_1_mult_513_C418_n222), .D(dp_cluster_1_mult_513_C418_n219), 
        .CO(dp_cluster_1_mult_513_C418_n216), .COX(
        dp_cluster_1_mult_513_C418_n215), .S(dp_cluster_1_mult_513_C418_n217)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U131 ( .A(
        dp_cluster_1_mult_513_C418_n324), .B(dp_cluster_1_mult_513_C418_n295), 
        .C(dp_cluster_1_mult_513_C418_n309), .CIX(
        dp_cluster_1_mult_513_C418_n220), .D(dp_cluster_1_mult_513_C418_n338), 
        .CO(dp_cluster_1_mult_513_C418_n213), .COX(
        dp_cluster_1_mult_513_C418_n212), .S(dp_cluster_1_mult_513_C418_n214)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U130 ( .A(
        dp_cluster_1_mult_513_C418_n352), .B(dp_cluster_1_mult_513_C418_n367), 
        .C(dp_cluster_1_mult_513_C418_n218), .CIX(
        dp_cluster_1_mult_513_C418_n214), .D(dp_cluster_1_mult_513_C418_n215), 
        .CO(dp_cluster_1_mult_513_C418_n210), .COX(
        dp_cluster_1_mult_513_C418_n209), .S(dp_cluster_1_mult_513_C418_n211)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U128 ( .A(
        dp_cluster_1_mult_513_C418_n366), .B(dp_cluster_1_mult_513_C418_n337), 
        .C(dp_cluster_1_mult_513_C418_n351), .CIX(
        dp_cluster_1_mult_513_C418_n212), .D(dp_cluster_1_mult_513_C418_n308), 
        .CO(dp_cluster_1_mult_513_C418_n205), .COX(
        dp_cluster_1_mult_513_C418_n204), .S(dp_cluster_1_mult_513_C418_n206)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U127 ( .A(
        dp_cluster_1_mult_513_C418_n208), .B(dp_cluster_1_mult_513_C418_n323), 
        .C(dp_cluster_1_mult_513_C418_n209), .CIX(
        dp_cluster_1_mult_513_C418_n213), .D(dp_cluster_1_mult_513_C418_n206), 
        .CO(dp_cluster_1_mult_513_C418_n202), .COX(
        dp_cluster_1_mult_513_C418_n201), .S(dp_cluster_1_mult_513_C418_n203)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U125 ( .A(
        dp_cluster_1_mult_513_C418_n322), .B(dp_cluster_1_mult_513_C418_n365), 
        .C(dp_cluster_1_mult_513_C418_n350), .CIX(
        dp_cluster_1_mult_513_C418_n200), .D(dp_cluster_1_mult_513_C418_n207), 
        .CO(dp_cluster_1_mult_513_C418_n197), .COX(
        dp_cluster_1_mult_513_C418_n196), .S(dp_cluster_1_mult_513_C418_n198)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U124 ( .A(
        dp_cluster_1_mult_513_C418_n204), .B(dp_cluster_1_mult_513_C418_n336), 
        .C(dp_cluster_1_mult_513_C418_n198), .CIX(
        dp_cluster_1_mult_513_C418_n201), .D(dp_cluster_1_mult_513_C418_n205), 
        .CO(dp_cluster_1_mult_513_C418_n194), .COX(
        dp_cluster_1_mult_513_C418_n193), .S(dp_cluster_1_mult_513_C418_n195)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U121 ( .A(
        dp_cluster_1_mult_513_C418_n306), .B(dp_cluster_1_mult_513_C418_n349), 
        .C(dp_cluster_1_mult_513_C418_n335), .CIX(
        dp_cluster_1_mult_513_C418_n190), .D(dp_cluster_1_mult_513_C418_n192), 
        .CO(dp_cluster_1_mult_513_C418_n187), .COX(
        dp_cluster_1_mult_513_C418_n186), .S(dp_cluster_1_mult_513_C418_n188)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U120 ( .A(
        dp_cluster_1_mult_513_C418_n199), .B(dp_cluster_1_mult_513_C418_n196), 
        .C(dp_cluster_1_mult_513_C418_n188), .CIX(
        dp_cluster_1_mult_513_C418_n193), .D(dp_cluster_1_mult_513_C418_n197), 
        .CO(dp_cluster_1_mult_513_C418_n184), .COX(
        dp_cluster_1_mult_513_C418_n183), .S(dp_cluster_1_mult_513_C418_n185)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U119 ( .A(
        dp_cluster_1_mult_513_C418_n291), .B(dp_cluster_1_mult_513_C418_n264), 
        .C(dp_cluster_1_mult_513_C418_n278), .CIX(
        dp_cluster_1_mult_513_C418_n191), .D(dp_cluster_1_mult_513_C418_n305), 
        .CO(dp_cluster_1_mult_513_C418_n181), .COX(
        dp_cluster_1_mult_513_C418_n180), .S(dp_cluster_1_mult_513_C418_n182)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U118 ( .A(
        dp_cluster_1_mult_513_C418_n363), .B(dp_cluster_1_mult_513_C418_n334), 
        .C(dp_cluster_1_mult_513_C418_n348), .CIX(
        dp_cluster_1_mult_513_C418_n189), .D(dp_cluster_1_mult_513_C418_n320), 
        .CO(dp_cluster_1_mult_513_C418_n178), .COX(
        dp_cluster_1_mult_513_C418_n177), .S(dp_cluster_1_mult_513_C418_n179)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U117 ( .A(
        dp_cluster_1_mult_513_C418_n182), .B(dp_cluster_1_mult_513_C418_n186), 
        .C(dp_cluster_1_mult_513_C418_n179), .CIX(
        dp_cluster_1_mult_513_C418_n183), .D(dp_cluster_1_mult_513_C418_n187), 
        .CO(dp_cluster_1_mult_513_C418_n175), .COX(
        dp_cluster_1_mult_513_C418_n174), .S(dp_cluster_1_mult_513_C418_n176)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U115 ( .A(
        dp_cluster_1_mult_513_C418_n362), .B(dp_cluster_1_mult_513_C418_n304), 
        .C(dp_cluster_1_mult_513_C418_n347), .CIX(
        dp_cluster_1_mult_513_C418_n180), .D(dp_cluster_1_mult_513_C418_n333), 
        .CO(dp_cluster_1_mult_513_C418_n170), .COX(
        dp_cluster_1_mult_513_C418_n169), .S(dp_cluster_1_mult_513_C418_n171)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U114 ( .A(
        dp_cluster_1_mult_513_C418_n277), .B(dp_cluster_1_mult_513_C418_n319), 
        .C(dp_cluster_1_mult_513_C418_n290), .CIX(
        dp_cluster_1_mult_513_C418_n177), .D(dp_cluster_1_mult_513_C418_n173), 
        .CO(dp_cluster_1_mult_513_C418_n167), .COX(
        dp_cluster_1_mult_513_C418_n166), .S(dp_cluster_1_mult_513_C418_n168)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U113 ( .A(
        dp_cluster_1_mult_513_C418_n168), .B(dp_cluster_1_mult_513_C418_n171), 
        .C(dp_cluster_1_mult_513_C418_n178), .CIX(
        dp_cluster_1_mult_513_C418_n174), .D(dp_cluster_1_mult_513_C418_n181), 
        .CO(dp_cluster_1_mult_513_C418_n164), .COX(
        dp_cluster_1_mult_513_C418_n163), .S(dp_cluster_1_mult_513_C418_n165)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U110 ( .A(
        dp_cluster_1_mult_513_C418_n262), .B(dp_cluster_1_mult_513_C418_n289), 
        .C(dp_cluster_1_mult_513_C418_n361), .CIX(
        dp_cluster_1_mult_513_C418_n169), .D(dp_cluster_1_mult_513_C418_n172), 
        .CO(dp_cluster_1_mult_513_C418_n159), .COX(
        dp_cluster_1_mult_513_C418_n158), .S(dp_cluster_1_mult_513_C418_n160)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U109 ( .A(
        dp_cluster_1_mult_513_C418_n303), .B(dp_cluster_1_mult_513_C418_n346), 
        .C(dp_cluster_1_mult_513_C418_n332), .CIX(
        dp_cluster_1_mult_513_C418_n166), .D(dp_cluster_1_mult_513_C418_n162), 
        .CO(dp_cluster_1_mult_513_C418_n156), .COX(
        dp_cluster_1_mult_513_C418_n155), .S(dp_cluster_1_mult_513_C418_n157)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U108 ( .A(
        dp_cluster_1_mult_513_C418_n170), .B(dp_cluster_1_mult_513_C418_n160), 
        .C(dp_cluster_1_mult_513_C418_n167), .CIX(
        dp_cluster_1_mult_513_C418_n163), .D(dp_cluster_1_mult_513_C418_n157), 
        .CO(dp_cluster_1_mult_513_C418_n153), .COX(
        dp_cluster_1_mult_513_C418_n152), .S(dp_cluster_1_mult_513_C418_n154)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U106 ( .A(
        dp_cluster_1_mult_513_C418_n331), .B(dp_cluster_1_mult_513_C418_n275), 
        .C(n1303), .CIX(dp_cluster_1_mult_513_C418_n158), .D(
        dp_cluster_1_mult_513_C418_n161), .CO(dp_cluster_1_mult_513_C418_n148), 
        .COX(dp_cluster_1_mult_513_C418_n147), .S(
        dp_cluster_1_mult_513_C418_n149) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U105 ( .A(
        dp_cluster_1_mult_513_C418_n317), .B(dp_cluster_1_mult_513_C418_n288), 
        .C(dp_cluster_1_mult_513_C418_n302), .CIX(
        dp_cluster_1_mult_513_C418_n155), .D(dp_cluster_1_mult_513_C418_n261), 
        .CO(dp_cluster_1_mult_513_C418_n145), .COX(
        dp_cluster_1_mult_513_C418_n144), .S(dp_cluster_1_mult_513_C418_n146)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U104 ( .A(
        dp_cluster_1_mult_513_C418_n149), .B(dp_cluster_1_mult_513_C418_n146), 
        .C(dp_cluster_1_mult_513_C418_n156), .CIX(
        dp_cluster_1_mult_513_C418_n152), .D(dp_cluster_1_mult_513_C418_n159), 
        .CO(dp_cluster_1_mult_513_C418_n142), .COX(
        dp_cluster_1_mult_513_C418_n141), .S(dp_cluster_1_mult_513_C418_n143)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U103 ( .A(
        dp_cluster_1_mult_513_C418_n150), .B(dp_cluster_1_mult_513_C418_n260), 
        .C(dp_cluster_1_mult_513_C418_n274), .CIX(
        dp_cluster_1_mult_513_C418_n147), .D(dp_cluster_1_mult_513_C418_n345), 
        .CO(dp_cluster_1_mult_513_C418_n139), .COX(
        dp_cluster_1_mult_513_C418_n138), .S(dp_cluster_1_mult_513_C418_n140)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U102 ( .A(
        dp_cluster_1_mult_513_C418_n330), .B(dp_cluster_1_mult_513_C418_n301), 
        .C(dp_cluster_1_mult_513_C418_n316), .CIX(
        dp_cluster_1_mult_513_C418_n144), .D(dp_cluster_1_mult_513_C418_n287), 
        .CO(dp_cluster_1_mult_513_C418_n136), .COX(
        dp_cluster_1_mult_513_C418_n135), .S(dp_cluster_1_mult_513_C418_n137)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U101 ( .A(
        dp_cluster_1_mult_513_C418_n140), .B(dp_cluster_1_mult_513_C418_n137), 
        .C(dp_cluster_1_mult_513_C418_n145), .CIX(
        dp_cluster_1_mult_513_C418_n141), .D(dp_cluster_1_mult_513_C418_n148), 
        .CO(dp_cluster_1_mult_513_C418_n133), .COX(
        dp_cluster_1_mult_513_C418_n132), .S(dp_cluster_1_mult_513_C418_n134)
         );
  CMPE42D1 dp_cluster_1_mult_513_C418_U98 ( .A(dp_cluster_1_mult_513_C418_n259), .B(dp_cluster_1_mult_513_C418_n300), .C(dp_cluster_1_mult_513_C418_n286), 
        .CIX(dp_cluster_1_mult_513_C418_n129), .D(
        dp_cluster_1_mult_513_C418_n135), .CO(dp_cluster_1_mult_513_C418_n126), 
        .COX(dp_cluster_1_mult_513_C418_n125), .S(
        dp_cluster_1_mult_513_C418_n127) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U97 ( .A(dp_cluster_1_mult_513_C418_n139), .B(dp_cluster_1_mult_513_C418_n138), .C(dp_cluster_1_mult_513_C418_n136), 
        .CIX(dp_cluster_1_mult_513_C418_n132), .D(
        dp_cluster_1_mult_513_C418_n127), .CO(dp_cluster_1_mult_513_C418_n123), 
        .COX(dp_cluster_1_mult_513_C418_n122), .S(
        dp_cluster_1_mult_513_C418_n124) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U95 ( .A(dp_cluster_1_mult_513_C418_n314), .B(dp_cluster_1_mult_513_C418_n285), .C(dp_cluster_1_mult_513_C418_n299), 
        .CIX(dp_cluster_1_mult_513_C418_n121), .D(
        dp_cluster_1_mult_513_C418_n272), .CO(dp_cluster_1_mult_513_C418_n118), 
        .COX(dp_cluster_1_mult_513_C418_n117), .S(
        dp_cluster_1_mult_513_C418_n119) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U94 ( .A(dp_cluster_1_mult_513_C418_n128), .B(dp_cluster_1_mult_513_C418_n125), .C(dp_cluster_1_mult_513_C418_n119), 
        .CIX(dp_cluster_1_mult_513_C418_n122), .D(
        dp_cluster_1_mult_513_C418_n126), .CO(dp_cluster_1_mult_513_C418_n115), 
        .COX(dp_cluster_1_mult_513_C418_n114), .S(
        dp_cluster_1_mult_513_C418_n116) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U92 ( .A(dp_cluster_1_mult_513_C418_n313), .B(dp_cluster_1_mult_513_C418_n271), .C(dp_cluster_1_mult_513_C418_n298), 
        .CIX(dp_cluster_1_mult_513_C418_n120), .D(n1292), .CO(
        dp_cluster_1_mult_513_C418_n110), .COX(dp_cluster_1_mult_513_C418_n109), .S(dp_cluster_1_mult_513_C418_n111) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U91 ( .A(dp_cluster_1_mult_513_C418_n117), .B(dp_cluster_1_mult_513_C418_n257), .C(dp_cluster_1_mult_513_C418_n111), 
        .CIX(dp_cluster_1_mult_513_C418_n114), .D(
        dp_cluster_1_mult_513_C418_n118), .CO(dp_cluster_1_mult_513_C418_n107), 
        .COX(dp_cluster_1_mult_513_C418_n106), .S(
        dp_cluster_1_mult_513_C418_n108) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U90 ( .A(dp_cluster_1_mult_513_C418_n297), .B(dp_cluster_1_mult_513_C418_n256), .C(dp_cluster_1_mult_513_C418_n284), 
        .CIX(dp_cluster_1_mult_513_C418_n109), .D(
        dp_cluster_1_mult_513_C418_n312), .CO(dp_cluster_1_mult_513_C418_n104), 
        .COX(dp_cluster_1_mult_513_C418_n103), .S(
        dp_cluster_1_mult_513_C418_n105) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U89 ( .A(dp_cluster_1_mult_513_C418_n112), .B(dp_cluster_1_mult_513_C418_n270), .C(dp_cluster_1_mult_513_C418_n105), 
        .CIX(dp_cluster_1_mult_513_C418_n106), .D(
        dp_cluster_1_mult_513_C418_n110), .CO(dp_cluster_1_mult_513_C418_n101), 
        .COX(dp_cluster_1_mult_513_C418_n100), .S(
        dp_cluster_1_mult_513_C418_n102) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U86 ( .A(dp_cluster_1_mult_513_C418_n103), .B(dp_cluster_1_mult_513_C418_n283), .C(dp_cluster_1_mult_513_C418_n97), 
        .CIX(dp_cluster_1_mult_513_C418_n100), .D(
        dp_cluster_1_mult_513_C418_n104), .CO(dp_cluster_1_mult_513_C418_n94), 
        .COX(dp_cluster_1_mult_513_C418_n93), .S(
        dp_cluster_1_mult_513_C418_n95) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U84 ( .A(dp_cluster_1_mult_513_C418_n98), 
        .B(dp_cluster_1_mult_513_C418_n282), .C(dp_cluster_1_mult_513_C418_n96), .CIX(dp_cluster_1_mult_513_C418_n93), .D(dp_cluster_1_mult_513_C418_n92), 
        .CO(dp_cluster_1_mult_513_C418_n89), .COX(
        dp_cluster_1_mult_513_C418_n88), .S(dp_cluster_1_mult_513_C418_n90) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U82 ( .A(dp_cluster_1_mult_513_C418_n253), .B(dp_cluster_1_mult_513_C418_n267), .C(n1293), .CIX(
        dp_cluster_1_mult_513_C418_n88), .D(dp_cluster_1_mult_513_C418_n91), 
        .CO(dp_cluster_1_mult_513_C418_n84), .COX(
        dp_cluster_1_mult_513_C418_n83), .S(dp_cluster_1_mult_513_C418_n85) );
  CMPE42D1 dp_cluster_1_mult_513_C418_U81 ( .A(dp_cluster_1_mult_513_C418_n266), .B(dp_cluster_1_mult_513_C418_n86), .C(dp_cluster_1_mult_513_C418_n252), 
        .CIX(dp_cluster_1_mult_513_C418_n83), .D(
        dp_cluster_1_mult_513_C418_n281), .CO(dp_cluster_1_mult_513_C418_n81), 
        .COX(dp_cluster_1_mult_513_C418_n80), .S(
        dp_cluster_1_mult_513_C418_n82) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U139 ( .A(
        dp_cluster_0_mult_485_C412_n371), .B(dp_cluster_0_mult_485_C412_n328), 
        .C(dp_cluster_0_mult_485_C412_n342), .CIX(
        dp_cluster_0_mult_485_C412_n237), .D(dp_cluster_0_mult_485_C412_n356), 
        .CO(dp_cluster_0_mult_485_C412_n233), .COX(
        dp_cluster_0_mult_485_C412_n232), .S(dp_cluster_0_mult_485_C412_n234)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U137 ( .A(
        dp_cluster_0_mult_485_C412_n341), .B(dp_cluster_0_mult_485_C412_n370), 
        .C(dp_cluster_0_mult_485_C412_n355), .CIX(
        dp_cluster_0_mult_485_C412_n232), .D(dp_cluster_0_mult_485_C412_n231), 
        .CO(dp_cluster_0_mult_485_C412_n228), .COX(
        dp_cluster_0_mult_485_C412_n227), .S(dp_cluster_0_mult_485_C412_n229)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U135 ( .A(
        dp_cluster_0_mult_485_C412_n354), .B(dp_cluster_0_mult_485_C412_n369), 
        .C(dp_cluster_0_mult_485_C412_n230), .CIX(
        dp_cluster_0_mult_485_C412_n226), .D(dp_cluster_0_mult_485_C412_n227), 
        .CO(dp_cluster_0_mult_485_C412_n223), .COX(
        dp_cluster_0_mult_485_C412_n222), .S(dp_cluster_0_mult_485_C412_n224)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U132 ( .A(
        dp_cluster_0_mult_485_C412_n221), .B(dp_cluster_0_mult_485_C412_n368), 
        .C(dp_cluster_0_mult_485_C412_n225), .CIX(
        dp_cluster_0_mult_485_C412_n222), .D(dp_cluster_0_mult_485_C412_n219), 
        .CO(dp_cluster_0_mult_485_C412_n216), .COX(
        dp_cluster_0_mult_485_C412_n215), .S(dp_cluster_0_mult_485_C412_n217)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U131 ( .A(
        dp_cluster_0_mult_485_C412_n324), .B(dp_cluster_0_mult_485_C412_n295), 
        .C(dp_cluster_0_mult_485_C412_n309), .CIX(
        dp_cluster_0_mult_485_C412_n220), .D(dp_cluster_0_mult_485_C412_n338), 
        .CO(dp_cluster_0_mult_485_C412_n213), .COX(
        dp_cluster_0_mult_485_C412_n212), .S(dp_cluster_0_mult_485_C412_n214)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U130 ( .A(
        dp_cluster_0_mult_485_C412_n352), .B(dp_cluster_0_mult_485_C412_n367), 
        .C(dp_cluster_0_mult_485_C412_n218), .CIX(
        dp_cluster_0_mult_485_C412_n214), .D(dp_cluster_0_mult_485_C412_n215), 
        .CO(dp_cluster_0_mult_485_C412_n210), .COX(
        dp_cluster_0_mult_485_C412_n209), .S(dp_cluster_0_mult_485_C412_n211)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U128 ( .A(
        dp_cluster_0_mult_485_C412_n366), .B(dp_cluster_0_mult_485_C412_n337), 
        .C(dp_cluster_0_mult_485_C412_n351), .CIX(
        dp_cluster_0_mult_485_C412_n212), .D(dp_cluster_0_mult_485_C412_n308), 
        .CO(dp_cluster_0_mult_485_C412_n205), .COX(
        dp_cluster_0_mult_485_C412_n204), .S(dp_cluster_0_mult_485_C412_n206)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U127 ( .A(
        dp_cluster_0_mult_485_C412_n208), .B(dp_cluster_0_mult_485_C412_n323), 
        .C(dp_cluster_0_mult_485_C412_n209), .CIX(
        dp_cluster_0_mult_485_C412_n213), .D(dp_cluster_0_mult_485_C412_n206), 
        .CO(dp_cluster_0_mult_485_C412_n202), .COX(
        dp_cluster_0_mult_485_C412_n201), .S(dp_cluster_0_mult_485_C412_n203)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U125 ( .A(
        dp_cluster_0_mult_485_C412_n322), .B(dp_cluster_0_mult_485_C412_n365), 
        .C(dp_cluster_0_mult_485_C412_n350), .CIX(
        dp_cluster_0_mult_485_C412_n200), .D(dp_cluster_0_mult_485_C412_n207), 
        .CO(dp_cluster_0_mult_485_C412_n197), .COX(
        dp_cluster_0_mult_485_C412_n196), .S(dp_cluster_0_mult_485_C412_n198)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U124 ( .A(
        dp_cluster_0_mult_485_C412_n204), .B(dp_cluster_0_mult_485_C412_n336), 
        .C(dp_cluster_0_mult_485_C412_n198), .CIX(
        dp_cluster_0_mult_485_C412_n201), .D(dp_cluster_0_mult_485_C412_n205), 
        .CO(dp_cluster_0_mult_485_C412_n194), .COX(
        dp_cluster_0_mult_485_C412_n193), .S(dp_cluster_0_mult_485_C412_n195)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U121 ( .A(
        dp_cluster_0_mult_485_C412_n306), .B(dp_cluster_0_mult_485_C412_n349), 
        .C(dp_cluster_0_mult_485_C412_n335), .CIX(
        dp_cluster_0_mult_485_C412_n190), .D(dp_cluster_0_mult_485_C412_n192), 
        .CO(dp_cluster_0_mult_485_C412_n187), .COX(
        dp_cluster_0_mult_485_C412_n186), .S(dp_cluster_0_mult_485_C412_n188)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U120 ( .A(
        dp_cluster_0_mult_485_C412_n199), .B(dp_cluster_0_mult_485_C412_n196), 
        .C(dp_cluster_0_mult_485_C412_n188), .CIX(
        dp_cluster_0_mult_485_C412_n193), .D(dp_cluster_0_mult_485_C412_n197), 
        .CO(dp_cluster_0_mult_485_C412_n184), .COX(
        dp_cluster_0_mult_485_C412_n183), .S(dp_cluster_0_mult_485_C412_n185)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U119 ( .A(
        dp_cluster_0_mult_485_C412_n291), .B(dp_cluster_0_mult_485_C412_n264), 
        .C(dp_cluster_0_mult_485_C412_n278), .CIX(
        dp_cluster_0_mult_485_C412_n191), .D(dp_cluster_0_mult_485_C412_n305), 
        .CO(dp_cluster_0_mult_485_C412_n181), .COX(
        dp_cluster_0_mult_485_C412_n180), .S(dp_cluster_0_mult_485_C412_n182)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U118 ( .A(
        dp_cluster_0_mult_485_C412_n363), .B(dp_cluster_0_mult_485_C412_n334), 
        .C(dp_cluster_0_mult_485_C412_n348), .CIX(
        dp_cluster_0_mult_485_C412_n189), .D(dp_cluster_0_mult_485_C412_n320), 
        .CO(dp_cluster_0_mult_485_C412_n178), .COX(
        dp_cluster_0_mult_485_C412_n177), .S(dp_cluster_0_mult_485_C412_n179)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U117 ( .A(
        dp_cluster_0_mult_485_C412_n182), .B(dp_cluster_0_mult_485_C412_n186), 
        .C(dp_cluster_0_mult_485_C412_n179), .CIX(
        dp_cluster_0_mult_485_C412_n183), .D(dp_cluster_0_mult_485_C412_n187), 
        .CO(dp_cluster_0_mult_485_C412_n175), .COX(
        dp_cluster_0_mult_485_C412_n174), .S(dp_cluster_0_mult_485_C412_n176)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U115 ( .A(
        dp_cluster_0_mult_485_C412_n362), .B(dp_cluster_0_mult_485_C412_n304), 
        .C(dp_cluster_0_mult_485_C412_n347), .CIX(
        dp_cluster_0_mult_485_C412_n180), .D(dp_cluster_0_mult_485_C412_n333), 
        .CO(dp_cluster_0_mult_485_C412_n170), .COX(
        dp_cluster_0_mult_485_C412_n169), .S(dp_cluster_0_mult_485_C412_n171)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U114 ( .A(
        dp_cluster_0_mult_485_C412_n277), .B(dp_cluster_0_mult_485_C412_n319), 
        .C(dp_cluster_0_mult_485_C412_n290), .CIX(
        dp_cluster_0_mult_485_C412_n177), .D(dp_cluster_0_mult_485_C412_n173), 
        .CO(dp_cluster_0_mult_485_C412_n167), .COX(
        dp_cluster_0_mult_485_C412_n166), .S(dp_cluster_0_mult_485_C412_n168)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U113 ( .A(
        dp_cluster_0_mult_485_C412_n168), .B(dp_cluster_0_mult_485_C412_n171), 
        .C(dp_cluster_0_mult_485_C412_n178), .CIX(
        dp_cluster_0_mult_485_C412_n174), .D(dp_cluster_0_mult_485_C412_n181), 
        .CO(dp_cluster_0_mult_485_C412_n164), .COX(
        dp_cluster_0_mult_485_C412_n163), .S(dp_cluster_0_mult_485_C412_n165)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U110 ( .A(
        dp_cluster_0_mult_485_C412_n262), .B(dp_cluster_0_mult_485_C412_n289), 
        .C(dp_cluster_0_mult_485_C412_n361), .CIX(
        dp_cluster_0_mult_485_C412_n169), .D(dp_cluster_0_mult_485_C412_n172), 
        .CO(dp_cluster_0_mult_485_C412_n159), .COX(
        dp_cluster_0_mult_485_C412_n158), .S(dp_cluster_0_mult_485_C412_n160)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U109 ( .A(
        dp_cluster_0_mult_485_C412_n303), .B(dp_cluster_0_mult_485_C412_n346), 
        .C(dp_cluster_0_mult_485_C412_n332), .CIX(
        dp_cluster_0_mult_485_C412_n166), .D(dp_cluster_0_mult_485_C412_n162), 
        .CO(dp_cluster_0_mult_485_C412_n156), .COX(
        dp_cluster_0_mult_485_C412_n155), .S(dp_cluster_0_mult_485_C412_n157)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U108 ( .A(
        dp_cluster_0_mult_485_C412_n170), .B(dp_cluster_0_mult_485_C412_n160), 
        .C(dp_cluster_0_mult_485_C412_n167), .CIX(
        dp_cluster_0_mult_485_C412_n163), .D(dp_cluster_0_mult_485_C412_n157), 
        .CO(dp_cluster_0_mult_485_C412_n153), .COX(
        dp_cluster_0_mult_485_C412_n152), .S(dp_cluster_0_mult_485_C412_n154)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U106 ( .A(
        dp_cluster_0_mult_485_C412_n331), .B(dp_cluster_0_mult_485_C412_n275), 
        .C(n1170), .CIX(dp_cluster_0_mult_485_C412_n158), .D(
        dp_cluster_0_mult_485_C412_n161), .CO(dp_cluster_0_mult_485_C412_n148), 
        .COX(dp_cluster_0_mult_485_C412_n147), .S(
        dp_cluster_0_mult_485_C412_n149) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U105 ( .A(
        dp_cluster_0_mult_485_C412_n317), .B(dp_cluster_0_mult_485_C412_n288), 
        .C(dp_cluster_0_mult_485_C412_n302), .CIX(
        dp_cluster_0_mult_485_C412_n155), .D(dp_cluster_0_mult_485_C412_n261), 
        .CO(dp_cluster_0_mult_485_C412_n145), .COX(
        dp_cluster_0_mult_485_C412_n144), .S(dp_cluster_0_mult_485_C412_n146)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U104 ( .A(
        dp_cluster_0_mult_485_C412_n149), .B(dp_cluster_0_mult_485_C412_n146), 
        .C(dp_cluster_0_mult_485_C412_n156), .CIX(
        dp_cluster_0_mult_485_C412_n152), .D(dp_cluster_0_mult_485_C412_n159), 
        .CO(dp_cluster_0_mult_485_C412_n142), .COX(
        dp_cluster_0_mult_485_C412_n141), .S(dp_cluster_0_mult_485_C412_n143)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U103 ( .A(
        dp_cluster_0_mult_485_C412_n150), .B(dp_cluster_0_mult_485_C412_n260), 
        .C(dp_cluster_0_mult_485_C412_n274), .CIX(
        dp_cluster_0_mult_485_C412_n147), .D(dp_cluster_0_mult_485_C412_n345), 
        .CO(dp_cluster_0_mult_485_C412_n139), .COX(
        dp_cluster_0_mult_485_C412_n138), .S(dp_cluster_0_mult_485_C412_n140)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U102 ( .A(
        dp_cluster_0_mult_485_C412_n330), .B(dp_cluster_0_mult_485_C412_n301), 
        .C(dp_cluster_0_mult_485_C412_n316), .CIX(
        dp_cluster_0_mult_485_C412_n144), .D(dp_cluster_0_mult_485_C412_n287), 
        .CO(dp_cluster_0_mult_485_C412_n136), .COX(
        dp_cluster_0_mult_485_C412_n135), .S(dp_cluster_0_mult_485_C412_n137)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U101 ( .A(
        dp_cluster_0_mult_485_C412_n140), .B(dp_cluster_0_mult_485_C412_n137), 
        .C(dp_cluster_0_mult_485_C412_n145), .CIX(
        dp_cluster_0_mult_485_C412_n141), .D(dp_cluster_0_mult_485_C412_n148), 
        .CO(dp_cluster_0_mult_485_C412_n133), .COX(
        dp_cluster_0_mult_485_C412_n132), .S(dp_cluster_0_mult_485_C412_n134)
         );
  CMPE42D1 dp_cluster_0_mult_485_C412_U98 ( .A(dp_cluster_0_mult_485_C412_n259), .B(dp_cluster_0_mult_485_C412_n300), .C(dp_cluster_0_mult_485_C412_n286), 
        .CIX(dp_cluster_0_mult_485_C412_n129), .D(
        dp_cluster_0_mult_485_C412_n135), .CO(dp_cluster_0_mult_485_C412_n126), 
        .COX(dp_cluster_0_mult_485_C412_n125), .S(
        dp_cluster_0_mult_485_C412_n127) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U97 ( .A(dp_cluster_0_mult_485_C412_n139), .B(dp_cluster_0_mult_485_C412_n138), .C(dp_cluster_0_mult_485_C412_n136), 
        .CIX(dp_cluster_0_mult_485_C412_n132), .D(
        dp_cluster_0_mult_485_C412_n127), .CO(dp_cluster_0_mult_485_C412_n123), 
        .COX(dp_cluster_0_mult_485_C412_n122), .S(
        dp_cluster_0_mult_485_C412_n124) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U95 ( .A(dp_cluster_0_mult_485_C412_n314), .B(dp_cluster_0_mult_485_C412_n285), .C(dp_cluster_0_mult_485_C412_n299), 
        .CIX(dp_cluster_0_mult_485_C412_n121), .D(
        dp_cluster_0_mult_485_C412_n272), .CO(dp_cluster_0_mult_485_C412_n118), 
        .COX(dp_cluster_0_mult_485_C412_n117), .S(
        dp_cluster_0_mult_485_C412_n119) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U94 ( .A(dp_cluster_0_mult_485_C412_n128), .B(dp_cluster_0_mult_485_C412_n125), .C(dp_cluster_0_mult_485_C412_n119), 
        .CIX(dp_cluster_0_mult_485_C412_n122), .D(
        dp_cluster_0_mult_485_C412_n126), .CO(dp_cluster_0_mult_485_C412_n115), 
        .COX(dp_cluster_0_mult_485_C412_n114), .S(
        dp_cluster_0_mult_485_C412_n116) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U92 ( .A(dp_cluster_0_mult_485_C412_n313), .B(dp_cluster_0_mult_485_C412_n271), .C(dp_cluster_0_mult_485_C412_n298), 
        .CIX(dp_cluster_0_mult_485_C412_n120), .D(n1154), .CO(
        dp_cluster_0_mult_485_C412_n110), .COX(dp_cluster_0_mult_485_C412_n109), .S(dp_cluster_0_mult_485_C412_n111) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U91 ( .A(dp_cluster_0_mult_485_C412_n117), .B(dp_cluster_0_mult_485_C412_n257), .C(dp_cluster_0_mult_485_C412_n111), 
        .CIX(dp_cluster_0_mult_485_C412_n114), .D(
        dp_cluster_0_mult_485_C412_n118), .CO(dp_cluster_0_mult_485_C412_n107), 
        .COX(dp_cluster_0_mult_485_C412_n106), .S(
        dp_cluster_0_mult_485_C412_n108) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U90 ( .A(dp_cluster_0_mult_485_C412_n297), .B(dp_cluster_0_mult_485_C412_n256), .C(dp_cluster_0_mult_485_C412_n284), 
        .CIX(dp_cluster_0_mult_485_C412_n109), .D(
        dp_cluster_0_mult_485_C412_n312), .CO(dp_cluster_0_mult_485_C412_n104), 
        .COX(dp_cluster_0_mult_485_C412_n103), .S(
        dp_cluster_0_mult_485_C412_n105) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U89 ( .A(dp_cluster_0_mult_485_C412_n112), .B(dp_cluster_0_mult_485_C412_n270), .C(dp_cluster_0_mult_485_C412_n105), 
        .CIX(dp_cluster_0_mult_485_C412_n106), .D(
        dp_cluster_0_mult_485_C412_n110), .CO(dp_cluster_0_mult_485_C412_n101), 
        .COX(dp_cluster_0_mult_485_C412_n100), .S(
        dp_cluster_0_mult_485_C412_n102) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U86 ( .A(dp_cluster_0_mult_485_C412_n103), .B(dp_cluster_0_mult_485_C412_n283), .C(dp_cluster_0_mult_485_C412_n97), 
        .CIX(dp_cluster_0_mult_485_C412_n100), .D(
        dp_cluster_0_mult_485_C412_n104), .CO(dp_cluster_0_mult_485_C412_n94), 
        .COX(dp_cluster_0_mult_485_C412_n93), .S(
        dp_cluster_0_mult_485_C412_n95) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U84 ( .A(dp_cluster_0_mult_485_C412_n98), 
        .B(dp_cluster_0_mult_485_C412_n282), .C(dp_cluster_0_mult_485_C412_n96), .CIX(dp_cluster_0_mult_485_C412_n93), .D(dp_cluster_0_mult_485_C412_n92), 
        .CO(dp_cluster_0_mult_485_C412_n89), .COX(
        dp_cluster_0_mult_485_C412_n88), .S(dp_cluster_0_mult_485_C412_n90) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U82 ( .A(dp_cluster_0_mult_485_C412_n253), .B(dp_cluster_0_mult_485_C412_n267), .C(n1156), .CIX(
        dp_cluster_0_mult_485_C412_n88), .D(dp_cluster_0_mult_485_C412_n91), 
        .CO(dp_cluster_0_mult_485_C412_n84), .COX(
        dp_cluster_0_mult_485_C412_n83), .S(dp_cluster_0_mult_485_C412_n85) );
  CMPE42D1 dp_cluster_0_mult_485_C412_U81 ( .A(dp_cluster_0_mult_485_C412_n266), .B(dp_cluster_0_mult_485_C412_n86), .C(dp_cluster_0_mult_485_C412_n252), 
        .CIX(dp_cluster_0_mult_485_C412_n83), .D(
        dp_cluster_0_mult_485_C412_n281), .CO(dp_cluster_0_mult_485_C412_n81), 
        .COX(dp_cluster_0_mult_485_C412_n80), .S(
        dp_cluster_0_mult_485_C412_n82) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U139 ( .A(
        dp_cluster_0_mult_486_C412_n371), .B(dp_cluster_0_mult_486_C412_n328), 
        .C(dp_cluster_0_mult_486_C412_n342), .CIX(
        dp_cluster_0_mult_486_C412_n237), .D(dp_cluster_0_mult_486_C412_n356), 
        .CO(dp_cluster_0_mult_486_C412_n233), .COX(
        dp_cluster_0_mult_486_C412_n232), .S(dp_cluster_0_mult_486_C412_n234)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U137 ( .A(
        dp_cluster_0_mult_486_C412_n341), .B(dp_cluster_0_mult_486_C412_n370), 
        .C(dp_cluster_0_mult_486_C412_n355), .CIX(
        dp_cluster_0_mult_486_C412_n232), .D(dp_cluster_0_mult_486_C412_n231), 
        .CO(dp_cluster_0_mult_486_C412_n228), .COX(
        dp_cluster_0_mult_486_C412_n227), .S(dp_cluster_0_mult_486_C412_n229)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U135 ( .A(
        dp_cluster_0_mult_486_C412_n354), .B(dp_cluster_0_mult_486_C412_n369), 
        .C(dp_cluster_0_mult_486_C412_n230), .CIX(
        dp_cluster_0_mult_486_C412_n226), .D(dp_cluster_0_mult_486_C412_n227), 
        .CO(dp_cluster_0_mult_486_C412_n223), .COX(
        dp_cluster_0_mult_486_C412_n222), .S(dp_cluster_0_mult_486_C412_n224)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U132 ( .A(
        dp_cluster_0_mult_486_C412_n221), .B(dp_cluster_0_mult_486_C412_n368), 
        .C(dp_cluster_0_mult_486_C412_n225), .CIX(
        dp_cluster_0_mult_486_C412_n222), .D(dp_cluster_0_mult_486_C412_n219), 
        .CO(dp_cluster_0_mult_486_C412_n216), .COX(
        dp_cluster_0_mult_486_C412_n215), .S(dp_cluster_0_mult_486_C412_n217)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U131 ( .A(
        dp_cluster_0_mult_486_C412_n324), .B(dp_cluster_0_mult_486_C412_n295), 
        .C(dp_cluster_0_mult_486_C412_n309), .CIX(
        dp_cluster_0_mult_486_C412_n220), .D(dp_cluster_0_mult_486_C412_n338), 
        .CO(dp_cluster_0_mult_486_C412_n213), .COX(
        dp_cluster_0_mult_486_C412_n212), .S(dp_cluster_0_mult_486_C412_n214)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U130 ( .A(
        dp_cluster_0_mult_486_C412_n352), .B(dp_cluster_0_mult_486_C412_n367), 
        .C(dp_cluster_0_mult_486_C412_n218), .CIX(
        dp_cluster_0_mult_486_C412_n214), .D(dp_cluster_0_mult_486_C412_n215), 
        .CO(dp_cluster_0_mult_486_C412_n210), .COX(
        dp_cluster_0_mult_486_C412_n209), .S(dp_cluster_0_mult_486_C412_n211)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U128 ( .A(
        dp_cluster_0_mult_486_C412_n366), .B(dp_cluster_0_mult_486_C412_n337), 
        .C(dp_cluster_0_mult_486_C412_n351), .CIX(
        dp_cluster_0_mult_486_C412_n212), .D(dp_cluster_0_mult_486_C412_n308), 
        .CO(dp_cluster_0_mult_486_C412_n205), .COX(
        dp_cluster_0_mult_486_C412_n204), .S(dp_cluster_0_mult_486_C412_n206)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U127 ( .A(
        dp_cluster_0_mult_486_C412_n208), .B(dp_cluster_0_mult_486_C412_n323), 
        .C(dp_cluster_0_mult_486_C412_n209), .CIX(
        dp_cluster_0_mult_486_C412_n213), .D(dp_cluster_0_mult_486_C412_n206), 
        .CO(dp_cluster_0_mult_486_C412_n202), .COX(
        dp_cluster_0_mult_486_C412_n201), .S(dp_cluster_0_mult_486_C412_n203)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U125 ( .A(
        dp_cluster_0_mult_486_C412_n322), .B(dp_cluster_0_mult_486_C412_n365), 
        .C(dp_cluster_0_mult_486_C412_n350), .CIX(
        dp_cluster_0_mult_486_C412_n200), .D(dp_cluster_0_mult_486_C412_n207), 
        .CO(dp_cluster_0_mult_486_C412_n197), .COX(
        dp_cluster_0_mult_486_C412_n196), .S(dp_cluster_0_mult_486_C412_n198)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U124 ( .A(
        dp_cluster_0_mult_486_C412_n204), .B(dp_cluster_0_mult_486_C412_n336), 
        .C(dp_cluster_0_mult_486_C412_n198), .CIX(
        dp_cluster_0_mult_486_C412_n201), .D(dp_cluster_0_mult_486_C412_n205), 
        .CO(dp_cluster_0_mult_486_C412_n194), .COX(
        dp_cluster_0_mult_486_C412_n193), .S(dp_cluster_0_mult_486_C412_n195)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U121 ( .A(
        dp_cluster_0_mult_486_C412_n306), .B(dp_cluster_0_mult_486_C412_n349), 
        .C(dp_cluster_0_mult_486_C412_n335), .CIX(
        dp_cluster_0_mult_486_C412_n190), .D(dp_cluster_0_mult_486_C412_n192), 
        .CO(dp_cluster_0_mult_486_C412_n187), .COX(
        dp_cluster_0_mult_486_C412_n186), .S(dp_cluster_0_mult_486_C412_n188)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U120 ( .A(
        dp_cluster_0_mult_486_C412_n199), .B(dp_cluster_0_mult_486_C412_n196), 
        .C(dp_cluster_0_mult_486_C412_n188), .CIX(
        dp_cluster_0_mult_486_C412_n193), .D(dp_cluster_0_mult_486_C412_n197), 
        .CO(dp_cluster_0_mult_486_C412_n184), .COX(
        dp_cluster_0_mult_486_C412_n183), .S(dp_cluster_0_mult_486_C412_n185)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U119 ( .A(
        dp_cluster_0_mult_486_C412_n291), .B(dp_cluster_0_mult_486_C412_n264), 
        .C(dp_cluster_0_mult_486_C412_n278), .CIX(
        dp_cluster_0_mult_486_C412_n191), .D(dp_cluster_0_mult_486_C412_n305), 
        .CO(dp_cluster_0_mult_486_C412_n181), .COX(
        dp_cluster_0_mult_486_C412_n180), .S(dp_cluster_0_mult_486_C412_n182)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U118 ( .A(
        dp_cluster_0_mult_486_C412_n363), .B(dp_cluster_0_mult_486_C412_n334), 
        .C(dp_cluster_0_mult_486_C412_n348), .CIX(
        dp_cluster_0_mult_486_C412_n189), .D(dp_cluster_0_mult_486_C412_n320), 
        .CO(dp_cluster_0_mult_486_C412_n178), .COX(
        dp_cluster_0_mult_486_C412_n177), .S(dp_cluster_0_mult_486_C412_n179)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U117 ( .A(
        dp_cluster_0_mult_486_C412_n182), .B(dp_cluster_0_mult_486_C412_n186), 
        .C(dp_cluster_0_mult_486_C412_n179), .CIX(
        dp_cluster_0_mult_486_C412_n183), .D(dp_cluster_0_mult_486_C412_n187), 
        .CO(dp_cluster_0_mult_486_C412_n175), .COX(
        dp_cluster_0_mult_486_C412_n174), .S(dp_cluster_0_mult_486_C412_n176)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U115 ( .A(
        dp_cluster_0_mult_486_C412_n362), .B(dp_cluster_0_mult_486_C412_n304), 
        .C(dp_cluster_0_mult_486_C412_n347), .CIX(
        dp_cluster_0_mult_486_C412_n180), .D(dp_cluster_0_mult_486_C412_n333), 
        .CO(dp_cluster_0_mult_486_C412_n170), .COX(
        dp_cluster_0_mult_486_C412_n169), .S(dp_cluster_0_mult_486_C412_n171)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U114 ( .A(
        dp_cluster_0_mult_486_C412_n277), .B(dp_cluster_0_mult_486_C412_n319), 
        .C(dp_cluster_0_mult_486_C412_n290), .CIX(
        dp_cluster_0_mult_486_C412_n177), .D(dp_cluster_0_mult_486_C412_n173), 
        .CO(dp_cluster_0_mult_486_C412_n167), .COX(
        dp_cluster_0_mult_486_C412_n166), .S(dp_cluster_0_mult_486_C412_n168)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U113 ( .A(
        dp_cluster_0_mult_486_C412_n168), .B(dp_cluster_0_mult_486_C412_n171), 
        .C(dp_cluster_0_mult_486_C412_n178), .CIX(
        dp_cluster_0_mult_486_C412_n174), .D(dp_cluster_0_mult_486_C412_n181), 
        .CO(dp_cluster_0_mult_486_C412_n164), .COX(
        dp_cluster_0_mult_486_C412_n163), .S(dp_cluster_0_mult_486_C412_n165)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U110 ( .A(
        dp_cluster_0_mult_486_C412_n262), .B(dp_cluster_0_mult_486_C412_n289), 
        .C(dp_cluster_0_mult_486_C412_n361), .CIX(
        dp_cluster_0_mult_486_C412_n169), .D(dp_cluster_0_mult_486_C412_n172), 
        .CO(dp_cluster_0_mult_486_C412_n159), .COX(
        dp_cluster_0_mult_486_C412_n158), .S(dp_cluster_0_mult_486_C412_n160)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U109 ( .A(
        dp_cluster_0_mult_486_C412_n303), .B(dp_cluster_0_mult_486_C412_n346), 
        .C(dp_cluster_0_mult_486_C412_n332), .CIX(
        dp_cluster_0_mult_486_C412_n166), .D(dp_cluster_0_mult_486_C412_n162), 
        .CO(dp_cluster_0_mult_486_C412_n156), .COX(
        dp_cluster_0_mult_486_C412_n155), .S(dp_cluster_0_mult_486_C412_n157)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U108 ( .A(
        dp_cluster_0_mult_486_C412_n170), .B(dp_cluster_0_mult_486_C412_n160), 
        .C(dp_cluster_0_mult_486_C412_n167), .CIX(
        dp_cluster_0_mult_486_C412_n163), .D(dp_cluster_0_mult_486_C412_n157), 
        .CO(dp_cluster_0_mult_486_C412_n153), .COX(
        dp_cluster_0_mult_486_C412_n152), .S(dp_cluster_0_mult_486_C412_n154)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U106 ( .A(
        dp_cluster_0_mult_486_C412_n331), .B(dp_cluster_0_mult_486_C412_n275), 
        .C(n1302), .CIX(dp_cluster_0_mult_486_C412_n158), .D(
        dp_cluster_0_mult_486_C412_n161), .CO(dp_cluster_0_mult_486_C412_n148), 
        .COX(dp_cluster_0_mult_486_C412_n147), .S(
        dp_cluster_0_mult_486_C412_n149) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U105 ( .A(
        dp_cluster_0_mult_486_C412_n317), .B(dp_cluster_0_mult_486_C412_n288), 
        .C(dp_cluster_0_mult_486_C412_n302), .CIX(
        dp_cluster_0_mult_486_C412_n155), .D(dp_cluster_0_mult_486_C412_n261), 
        .CO(dp_cluster_0_mult_486_C412_n145), .COX(
        dp_cluster_0_mult_486_C412_n144), .S(dp_cluster_0_mult_486_C412_n146)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U104 ( .A(
        dp_cluster_0_mult_486_C412_n149), .B(dp_cluster_0_mult_486_C412_n146), 
        .C(dp_cluster_0_mult_486_C412_n156), .CIX(
        dp_cluster_0_mult_486_C412_n152), .D(dp_cluster_0_mult_486_C412_n159), 
        .CO(dp_cluster_0_mult_486_C412_n142), .COX(
        dp_cluster_0_mult_486_C412_n141), .S(dp_cluster_0_mult_486_C412_n143)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U103 ( .A(
        dp_cluster_0_mult_486_C412_n150), .B(dp_cluster_0_mult_486_C412_n260), 
        .C(dp_cluster_0_mult_486_C412_n274), .CIX(
        dp_cluster_0_mult_486_C412_n147), .D(dp_cluster_0_mult_486_C412_n345), 
        .CO(dp_cluster_0_mult_486_C412_n139), .COX(
        dp_cluster_0_mult_486_C412_n138), .S(dp_cluster_0_mult_486_C412_n140)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U102 ( .A(
        dp_cluster_0_mult_486_C412_n330), .B(dp_cluster_0_mult_486_C412_n301), 
        .C(dp_cluster_0_mult_486_C412_n316), .CIX(
        dp_cluster_0_mult_486_C412_n144), .D(dp_cluster_0_mult_486_C412_n287), 
        .CO(dp_cluster_0_mult_486_C412_n136), .COX(
        dp_cluster_0_mult_486_C412_n135), .S(dp_cluster_0_mult_486_C412_n137)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U101 ( .A(
        dp_cluster_0_mult_486_C412_n140), .B(dp_cluster_0_mult_486_C412_n137), 
        .C(dp_cluster_0_mult_486_C412_n145), .CIX(
        dp_cluster_0_mult_486_C412_n141), .D(dp_cluster_0_mult_486_C412_n148), 
        .CO(dp_cluster_0_mult_486_C412_n133), .COX(
        dp_cluster_0_mult_486_C412_n132), .S(dp_cluster_0_mult_486_C412_n134)
         );
  CMPE42D1 dp_cluster_0_mult_486_C412_U98 ( .A(dp_cluster_0_mult_486_C412_n259), .B(dp_cluster_0_mult_486_C412_n300), .C(dp_cluster_0_mult_486_C412_n286), 
        .CIX(dp_cluster_0_mult_486_C412_n129), .D(
        dp_cluster_0_mult_486_C412_n135), .CO(dp_cluster_0_mult_486_C412_n126), 
        .COX(dp_cluster_0_mult_486_C412_n125), .S(
        dp_cluster_0_mult_486_C412_n127) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U97 ( .A(dp_cluster_0_mult_486_C412_n139), .B(dp_cluster_0_mult_486_C412_n138), .C(dp_cluster_0_mult_486_C412_n136), 
        .CIX(dp_cluster_0_mult_486_C412_n132), .D(
        dp_cluster_0_mult_486_C412_n127), .CO(dp_cluster_0_mult_486_C412_n123), 
        .COX(dp_cluster_0_mult_486_C412_n122), .S(
        dp_cluster_0_mult_486_C412_n124) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U95 ( .A(dp_cluster_0_mult_486_C412_n314), .B(dp_cluster_0_mult_486_C412_n285), .C(dp_cluster_0_mult_486_C412_n299), 
        .CIX(dp_cluster_0_mult_486_C412_n121), .D(
        dp_cluster_0_mult_486_C412_n272), .CO(dp_cluster_0_mult_486_C412_n118), 
        .COX(dp_cluster_0_mult_486_C412_n117), .S(
        dp_cluster_0_mult_486_C412_n119) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U94 ( .A(dp_cluster_0_mult_486_C412_n128), .B(dp_cluster_0_mult_486_C412_n125), .C(dp_cluster_0_mult_486_C412_n119), 
        .CIX(dp_cluster_0_mult_486_C412_n122), .D(
        dp_cluster_0_mult_486_C412_n126), .CO(dp_cluster_0_mult_486_C412_n115), 
        .COX(dp_cluster_0_mult_486_C412_n114), .S(
        dp_cluster_0_mult_486_C412_n116) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U92 ( .A(dp_cluster_0_mult_486_C412_n313), .B(dp_cluster_0_mult_486_C412_n271), .C(dp_cluster_0_mult_486_C412_n298), 
        .CIX(dp_cluster_0_mult_486_C412_n120), .D(n1290), .CO(
        dp_cluster_0_mult_486_C412_n110), .COX(dp_cluster_0_mult_486_C412_n109), .S(dp_cluster_0_mult_486_C412_n111) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U91 ( .A(dp_cluster_0_mult_486_C412_n117), .B(dp_cluster_0_mult_486_C412_n257), .C(dp_cluster_0_mult_486_C412_n111), 
        .CIX(dp_cluster_0_mult_486_C412_n114), .D(
        dp_cluster_0_mult_486_C412_n118), .CO(dp_cluster_0_mult_486_C412_n107), 
        .COX(dp_cluster_0_mult_486_C412_n106), .S(
        dp_cluster_0_mult_486_C412_n108) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U90 ( .A(dp_cluster_0_mult_486_C412_n297), .B(dp_cluster_0_mult_486_C412_n256), .C(dp_cluster_0_mult_486_C412_n284), 
        .CIX(dp_cluster_0_mult_486_C412_n109), .D(
        dp_cluster_0_mult_486_C412_n312), .CO(dp_cluster_0_mult_486_C412_n104), 
        .COX(dp_cluster_0_mult_486_C412_n103), .S(
        dp_cluster_0_mult_486_C412_n105) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U89 ( .A(dp_cluster_0_mult_486_C412_n112), .B(dp_cluster_0_mult_486_C412_n270), .C(dp_cluster_0_mult_486_C412_n105), 
        .CIX(dp_cluster_0_mult_486_C412_n106), .D(
        dp_cluster_0_mult_486_C412_n110), .CO(dp_cluster_0_mult_486_C412_n101), 
        .COX(dp_cluster_0_mult_486_C412_n100), .S(
        dp_cluster_0_mult_486_C412_n102) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U86 ( .A(dp_cluster_0_mult_486_C412_n103), .B(dp_cluster_0_mult_486_C412_n283), .C(dp_cluster_0_mult_486_C412_n97), 
        .CIX(dp_cluster_0_mult_486_C412_n100), .D(
        dp_cluster_0_mult_486_C412_n104), .CO(dp_cluster_0_mult_486_C412_n94), 
        .COX(dp_cluster_0_mult_486_C412_n93), .S(
        dp_cluster_0_mult_486_C412_n95) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U84 ( .A(dp_cluster_0_mult_486_C412_n98), 
        .B(dp_cluster_0_mult_486_C412_n282), .C(dp_cluster_0_mult_486_C412_n96), .CIX(dp_cluster_0_mult_486_C412_n93), .D(dp_cluster_0_mult_486_C412_n92), 
        .CO(dp_cluster_0_mult_486_C412_n89), .COX(
        dp_cluster_0_mult_486_C412_n88), .S(dp_cluster_0_mult_486_C412_n90) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U82 ( .A(dp_cluster_0_mult_486_C412_n253), .B(dp_cluster_0_mult_486_C412_n267), .C(n1291), .CIX(
        dp_cluster_0_mult_486_C412_n88), .D(dp_cluster_0_mult_486_C412_n91), 
        .CO(dp_cluster_0_mult_486_C412_n84), .COX(
        dp_cluster_0_mult_486_C412_n83), .S(dp_cluster_0_mult_486_C412_n85) );
  CMPE42D1 dp_cluster_0_mult_486_C412_U81 ( .A(dp_cluster_0_mult_486_C412_n266), .B(dp_cluster_0_mult_486_C412_n86), .C(dp_cluster_0_mult_486_C412_n252), 
        .CIX(dp_cluster_0_mult_486_C412_n83), .D(
        dp_cluster_0_mult_486_C412_n281), .CO(dp_cluster_0_mult_486_C412_n81), 
        .COX(dp_cluster_0_mult_486_C412_n80), .S(
        dp_cluster_0_mult_486_C412_n82) );
  XOR3D1 add_328_U1_16 ( .A1(xi0_r[63]), .A2(xi4_r[63]), .A3(add_328_carry[16]), .Z(s1_0_r[16]) );
  XOR3D1 add_337_U1_16 ( .A1(xi0_i[63]), .A2(xi4_i[63]), .A3(add_337_carry[16]), .Z(s1_0_i[16]) );
  XOR3D1 add_329_U1_16 ( .A1(xi1_r[63]), .A2(xi5_r[63]), .A3(add_329_carry[16]), .Z(s1_1_r[16]) );
  XOR3D1 add_338_U1_16 ( .A1(xi1_i[63]), .A2(xi5_i[63]), .A3(add_338_carry[16]), .Z(s1_1_i[16]) );
  XOR3D1 add_330_U1_16 ( .A1(xi2_r[63]), .A2(xi6_r[63]), .A3(add_330_carry[16]), .Z(s1_2_r[16]) );
  XOR3D1 add_339_U1_16 ( .A1(xi2_i[63]), .A2(xi6_i[63]), .A3(add_339_carry[16]), .Z(s1_2_i[16]) );
  XOR3D1 add_331_U1_16 ( .A1(xi3_r[63]), .A2(xi7_r[63]), .A3(add_331_carry[16]), .Z(s1_3_r[16]) );
  XOR3D1 add_340_U1_16 ( .A1(xi3_i[63]), .A2(xi7_i[63]), .A3(add_340_carry[16]), .Z(s1_3_i[16]) );
  XOR3D1 sub_332_U2_16 ( .A1(xi0_r[63]), .A2(n1176), .A3(sub_332_carry[16]), 
        .Z(s1_4_r[16]) );
  XOR3D1 sub_341_U2_16 ( .A1(xi0_i[63]), .A2(n1306), .A3(sub_341_carry[16]), 
        .Z(s1_4_i[16]) );
  XOR3D1 sub_343_U2_16 ( .A1(xi2_i[63]), .A2(n1338), .A3(sub_343_carry[16]), 
        .Z(s1_6_i[16]) );
  XOR3D1 sub_334_U2_16 ( .A1(xi2_r[63]), .A2(n1208), .A3(sub_334_carry[16]), 
        .Z(s1_6_r[16]) );
  FA1D0 add_328_U1_15 ( .A(xi0_r[62]), .B(xi4_r[62]), .CI(add_328_carry[15]), 
        .CO(add_328_carry[16]), .S(s1_0_r[15]) );
  FA1D0 add_328_U1_14 ( .A(xi0_r[61]), .B(xi4_r[61]), .CI(add_328_carry[14]), 
        .CO(add_328_carry[15]), .S(s1_0_r[14]) );
  FA1D0 add_328_U1_13 ( .A(xi0_r[60]), .B(xi4_r[60]), .CI(add_328_carry[13]), 
        .CO(add_328_carry[14]), .S(s1_0_r[13]) );
  FA1D0 add_328_U1_12 ( .A(xi0_r[59]), .B(xi4_r[59]), .CI(add_328_carry[12]), 
        .CO(add_328_carry[13]), .S(s1_0_r[12]) );
  FA1D0 add_328_U1_11 ( .A(xi0_r[58]), .B(xi4_r[58]), .CI(add_328_carry[11]), 
        .CO(add_328_carry[12]), .S(s1_0_r[11]) );
  FA1D0 add_328_U1_10 ( .A(xi0_r[57]), .B(xi4_r[57]), .CI(add_328_carry[10]), 
        .CO(add_328_carry[11]), .S(s1_0_r[10]) );
  FA1D0 add_328_U1_9 ( .A(xi0_r[56]), .B(xi4_r[56]), .CI(add_328_carry[9]), 
        .CO(add_328_carry[10]), .S(s1_0_r[9]) );
  FA1D0 add_328_U1_8 ( .A(xi0_r[55]), .B(xi4_r[55]), .CI(add_328_carry[8]), 
        .CO(add_328_carry[9]), .S(s1_0_r[8]) );
  FA1D0 add_328_U1_7 ( .A(xi0_r[54]), .B(xi4_r[54]), .CI(add_328_carry[7]), 
        .CO(add_328_carry[8]), .S(s1_0_r[7]) );
  FA1D0 add_328_U1_6 ( .A(xi0_r[53]), .B(xi4_r[53]), .CI(add_328_carry[6]), 
        .CO(add_328_carry[7]), .S(s1_0_r[6]) );
  FA1D0 add_328_U1_5 ( .A(xi0_r[52]), .B(xi4_r[52]), .CI(add_328_carry[5]), 
        .CO(add_328_carry[6]), .S(s1_0_r[5]) );
  FA1D0 add_328_U1_4 ( .A(xi0_r[51]), .B(xi4_r[51]), .CI(add_328_carry[4]), 
        .CO(add_328_carry[5]), .S(s1_0_r[4]) );
  FA1D0 add_328_U1_3 ( .A(xi0_r[50]), .B(xi4_r[50]), .CI(add_328_carry[3]), 
        .CO(add_328_carry[4]), .S(s1_0_r[3]) );
  FA1D0 add_328_U1_2 ( .A(xi0_r[49]), .B(xi4_r[49]), .CI(add_328_carry[2]), 
        .CO(add_328_carry[3]), .S(s1_0_r[2]) );
  FA1D0 add_328_U1_1 ( .A(xi0_r[48]), .B(xi4_r[48]), .CI(add_328_carry[1]), 
        .CO(add_328_carry[2]), .S(s1_0_r[1]) );
  FA1D0 add_337_U1_15 ( .A(xi0_i[62]), .B(xi4_i[62]), .CI(add_337_carry[15]), 
        .CO(add_337_carry[16]), .S(s1_0_i[15]) );
  FA1D0 add_337_U1_14 ( .A(xi0_i[61]), .B(xi4_i[61]), .CI(add_337_carry[14]), 
        .CO(add_337_carry[15]), .S(s1_0_i[14]) );
  FA1D0 add_337_U1_13 ( .A(xi0_i[60]), .B(xi4_i[60]), .CI(add_337_carry[13]), 
        .CO(add_337_carry[14]), .S(s1_0_i[13]) );
  FA1D0 add_337_U1_12 ( .A(xi0_i[59]), .B(xi4_i[59]), .CI(add_337_carry[12]), 
        .CO(add_337_carry[13]), .S(s1_0_i[12]) );
  FA1D0 add_337_U1_11 ( .A(xi0_i[58]), .B(xi4_i[58]), .CI(add_337_carry[11]), 
        .CO(add_337_carry[12]), .S(s1_0_i[11]) );
  FA1D0 add_337_U1_10 ( .A(xi0_i[57]), .B(xi4_i[57]), .CI(add_337_carry[10]), 
        .CO(add_337_carry[11]), .S(s1_0_i[10]) );
  FA1D0 add_337_U1_9 ( .A(xi0_i[56]), .B(xi4_i[56]), .CI(add_337_carry[9]), 
        .CO(add_337_carry[10]), .S(s1_0_i[9]) );
  FA1D0 add_337_U1_8 ( .A(xi0_i[55]), .B(xi4_i[55]), .CI(add_337_carry[8]), 
        .CO(add_337_carry[9]), .S(s1_0_i[8]) );
  FA1D0 add_337_U1_7 ( .A(xi0_i[54]), .B(xi4_i[54]), .CI(add_337_carry[7]), 
        .CO(add_337_carry[8]), .S(s1_0_i[7]) );
  FA1D0 add_337_U1_6 ( .A(xi0_i[53]), .B(xi4_i[53]), .CI(add_337_carry[6]), 
        .CO(add_337_carry[7]), .S(s1_0_i[6]) );
  FA1D0 add_337_U1_5 ( .A(xi0_i[52]), .B(xi4_i[52]), .CI(add_337_carry[5]), 
        .CO(add_337_carry[6]), .S(s1_0_i[5]) );
  FA1D0 add_337_U1_4 ( .A(xi0_i[51]), .B(xi4_i[51]), .CI(add_337_carry[4]), 
        .CO(add_337_carry[5]), .S(s1_0_i[4]) );
  FA1D0 add_337_U1_3 ( .A(xi0_i[50]), .B(xi4_i[50]), .CI(add_337_carry[3]), 
        .CO(add_337_carry[4]), .S(s1_0_i[3]) );
  FA1D0 add_337_U1_2 ( .A(xi0_i[49]), .B(xi4_i[49]), .CI(add_337_carry[2]), 
        .CO(add_337_carry[3]), .S(s1_0_i[2]) );
  FA1D0 add_337_U1_1 ( .A(xi0_i[48]), .B(xi4_i[48]), .CI(add_337_carry[1]), 
        .CO(add_337_carry[2]), .S(s1_0_i[1]) );
  FA1D0 add_329_U1_15 ( .A(xi1_r[62]), .B(xi5_r[62]), .CI(add_329_carry[15]), 
        .CO(add_329_carry[16]), .S(s1_1_r[15]) );
  FA1D0 add_329_U1_14 ( .A(xi1_r[61]), .B(xi5_r[61]), .CI(add_329_carry[14]), 
        .CO(add_329_carry[15]), .S(s1_1_r[14]) );
  FA1D0 add_329_U1_13 ( .A(xi1_r[60]), .B(xi5_r[60]), .CI(add_329_carry[13]), 
        .CO(add_329_carry[14]), .S(s1_1_r[13]) );
  FA1D0 add_329_U1_12 ( .A(xi1_r[59]), .B(xi5_r[59]), .CI(add_329_carry[12]), 
        .CO(add_329_carry[13]), .S(s1_1_r[12]) );
  FA1D0 add_329_U1_11 ( .A(xi1_r[58]), .B(xi5_r[58]), .CI(add_329_carry[11]), 
        .CO(add_329_carry[12]), .S(s1_1_r[11]) );
  FA1D0 add_329_U1_10 ( .A(xi1_r[57]), .B(xi5_r[57]), .CI(add_329_carry[10]), 
        .CO(add_329_carry[11]), .S(s1_1_r[10]) );
  FA1D0 add_329_U1_9 ( .A(xi1_r[56]), .B(xi5_r[56]), .CI(add_329_carry[9]), 
        .CO(add_329_carry[10]), .S(s1_1_r[9]) );
  FA1D0 add_329_U1_8 ( .A(xi1_r[55]), .B(xi5_r[55]), .CI(add_329_carry[8]), 
        .CO(add_329_carry[9]), .S(s1_1_r[8]) );
  FA1D0 add_329_U1_7 ( .A(xi1_r[54]), .B(xi5_r[54]), .CI(add_329_carry[7]), 
        .CO(add_329_carry[8]), .S(s1_1_r[7]) );
  FA1D0 add_329_U1_6 ( .A(xi1_r[53]), .B(xi5_r[53]), .CI(add_329_carry[6]), 
        .CO(add_329_carry[7]), .S(s1_1_r[6]) );
  FA1D0 add_329_U1_5 ( .A(xi1_r[52]), .B(xi5_r[52]), .CI(add_329_carry[5]), 
        .CO(add_329_carry[6]), .S(s1_1_r[5]) );
  FA1D0 add_329_U1_4 ( .A(xi1_r[51]), .B(xi5_r[51]), .CI(add_329_carry[4]), 
        .CO(add_329_carry[5]), .S(s1_1_r[4]) );
  FA1D0 add_329_U1_3 ( .A(xi1_r[50]), .B(xi5_r[50]), .CI(add_329_carry[3]), 
        .CO(add_329_carry[4]), .S(s1_1_r[3]) );
  FA1D0 add_329_U1_2 ( .A(xi1_r[49]), .B(xi5_r[49]), .CI(add_329_carry[2]), 
        .CO(add_329_carry[3]), .S(s1_1_r[2]) );
  FA1D0 add_329_U1_1 ( .A(xi1_r[48]), .B(xi5_r[48]), .CI(add_329_carry[1]), 
        .CO(add_329_carry[2]), .S(s1_1_r[1]) );
  FA1D0 add_338_U1_15 ( .A(xi1_i[62]), .B(xi5_i[62]), .CI(add_338_carry[15]), 
        .CO(add_338_carry[16]), .S(s1_1_i[15]) );
  FA1D0 add_338_U1_14 ( .A(xi1_i[61]), .B(xi5_i[61]), .CI(add_338_carry[14]), 
        .CO(add_338_carry[15]), .S(s1_1_i[14]) );
  FA1D0 add_338_U1_13 ( .A(xi1_i[60]), .B(xi5_i[60]), .CI(add_338_carry[13]), 
        .CO(add_338_carry[14]), .S(s1_1_i[13]) );
  FA1D0 add_338_U1_12 ( .A(xi1_i[59]), .B(xi5_i[59]), .CI(add_338_carry[12]), 
        .CO(add_338_carry[13]), .S(s1_1_i[12]) );
  FA1D0 add_338_U1_11 ( .A(xi1_i[58]), .B(xi5_i[58]), .CI(add_338_carry[11]), 
        .CO(add_338_carry[12]), .S(s1_1_i[11]) );
  FA1D0 add_338_U1_10 ( .A(xi1_i[57]), .B(xi5_i[57]), .CI(add_338_carry[10]), 
        .CO(add_338_carry[11]), .S(s1_1_i[10]) );
  FA1D0 add_338_U1_9 ( .A(xi1_i[56]), .B(xi5_i[56]), .CI(add_338_carry[9]), 
        .CO(add_338_carry[10]), .S(s1_1_i[9]) );
  FA1D0 add_338_U1_8 ( .A(xi1_i[55]), .B(xi5_i[55]), .CI(add_338_carry[8]), 
        .CO(add_338_carry[9]), .S(s1_1_i[8]) );
  FA1D0 add_338_U1_7 ( .A(xi1_i[54]), .B(xi5_i[54]), .CI(add_338_carry[7]), 
        .CO(add_338_carry[8]), .S(s1_1_i[7]) );
  FA1D0 add_338_U1_6 ( .A(xi1_i[53]), .B(xi5_i[53]), .CI(add_338_carry[6]), 
        .CO(add_338_carry[7]), .S(s1_1_i[6]) );
  FA1D0 add_338_U1_5 ( .A(xi1_i[52]), .B(xi5_i[52]), .CI(add_338_carry[5]), 
        .CO(add_338_carry[6]), .S(s1_1_i[5]) );
  FA1D0 add_338_U1_4 ( .A(xi1_i[51]), .B(xi5_i[51]), .CI(add_338_carry[4]), 
        .CO(add_338_carry[5]), .S(s1_1_i[4]) );
  FA1D0 add_338_U1_3 ( .A(xi1_i[50]), .B(xi5_i[50]), .CI(add_338_carry[3]), 
        .CO(add_338_carry[4]), .S(s1_1_i[3]) );
  FA1D0 add_338_U1_2 ( .A(xi1_i[49]), .B(xi5_i[49]), .CI(add_338_carry[2]), 
        .CO(add_338_carry[3]), .S(s1_1_i[2]) );
  FA1D0 add_338_U1_1 ( .A(xi1_i[48]), .B(xi5_i[48]), .CI(add_338_carry[1]), 
        .CO(add_338_carry[2]), .S(s1_1_i[1]) );
  FA1D0 add_330_U1_15 ( .A(xi2_r[62]), .B(xi6_r[62]), .CI(add_330_carry[15]), 
        .CO(add_330_carry[16]), .S(s1_2_r[15]) );
  FA1D0 add_330_U1_14 ( .A(xi2_r[61]), .B(xi6_r[61]), .CI(add_330_carry[14]), 
        .CO(add_330_carry[15]), .S(s1_2_r[14]) );
  FA1D0 add_330_U1_13 ( .A(xi2_r[60]), .B(xi6_r[60]), .CI(add_330_carry[13]), 
        .CO(add_330_carry[14]), .S(s1_2_r[13]) );
  FA1D0 add_330_U1_12 ( .A(xi2_r[59]), .B(xi6_r[59]), .CI(add_330_carry[12]), 
        .CO(add_330_carry[13]), .S(s1_2_r[12]) );
  FA1D0 add_330_U1_11 ( .A(xi2_r[58]), .B(xi6_r[58]), .CI(add_330_carry[11]), 
        .CO(add_330_carry[12]), .S(s1_2_r[11]) );
  FA1D0 add_330_U1_10 ( .A(xi2_r[57]), .B(xi6_r[57]), .CI(add_330_carry[10]), 
        .CO(add_330_carry[11]), .S(s1_2_r[10]) );
  FA1D0 add_330_U1_9 ( .A(xi2_r[56]), .B(xi6_r[56]), .CI(add_330_carry[9]), 
        .CO(add_330_carry[10]), .S(s1_2_r[9]) );
  FA1D0 add_330_U1_8 ( .A(xi2_r[55]), .B(xi6_r[55]), .CI(add_330_carry[8]), 
        .CO(add_330_carry[9]), .S(s1_2_r[8]) );
  FA1D0 add_330_U1_7 ( .A(xi2_r[54]), .B(xi6_r[54]), .CI(add_330_carry[7]), 
        .CO(add_330_carry[8]), .S(s1_2_r[7]) );
  FA1D0 add_330_U1_6 ( .A(xi2_r[53]), .B(xi6_r[53]), .CI(add_330_carry[6]), 
        .CO(add_330_carry[7]), .S(s1_2_r[6]) );
  FA1D0 add_330_U1_5 ( .A(xi2_r[52]), .B(xi6_r[52]), .CI(add_330_carry[5]), 
        .CO(add_330_carry[6]), .S(s1_2_r[5]) );
  FA1D0 add_330_U1_4 ( .A(xi2_r[51]), .B(xi6_r[51]), .CI(add_330_carry[4]), 
        .CO(add_330_carry[5]), .S(s1_2_r[4]) );
  FA1D0 add_330_U1_3 ( .A(xi2_r[50]), .B(xi6_r[50]), .CI(add_330_carry[3]), 
        .CO(add_330_carry[4]), .S(s1_2_r[3]) );
  FA1D0 add_330_U1_2 ( .A(xi2_r[49]), .B(xi6_r[49]), .CI(add_330_carry[2]), 
        .CO(add_330_carry[3]), .S(s1_2_r[2]) );
  FA1D0 add_330_U1_1 ( .A(xi2_r[48]), .B(xi6_r[48]), .CI(add_330_carry[1]), 
        .CO(add_330_carry[2]), .S(s1_2_r[1]) );
  FA1D0 add_339_U1_15 ( .A(xi2_i[62]), .B(xi6_i[62]), .CI(add_339_carry[15]), 
        .CO(add_339_carry[16]), .S(s1_2_i[15]) );
  FA1D0 add_339_U1_14 ( .A(xi2_i[61]), .B(xi6_i[61]), .CI(add_339_carry[14]), 
        .CO(add_339_carry[15]), .S(s1_2_i[14]) );
  FA1D0 add_339_U1_13 ( .A(xi2_i[60]), .B(xi6_i[60]), .CI(add_339_carry[13]), 
        .CO(add_339_carry[14]), .S(s1_2_i[13]) );
  FA1D0 add_339_U1_12 ( .A(xi2_i[59]), .B(xi6_i[59]), .CI(add_339_carry[12]), 
        .CO(add_339_carry[13]), .S(s1_2_i[12]) );
  FA1D0 add_339_U1_11 ( .A(xi2_i[58]), .B(xi6_i[58]), .CI(add_339_carry[11]), 
        .CO(add_339_carry[12]), .S(s1_2_i[11]) );
  FA1D0 add_339_U1_10 ( .A(xi2_i[57]), .B(xi6_i[57]), .CI(add_339_carry[10]), 
        .CO(add_339_carry[11]), .S(s1_2_i[10]) );
  FA1D0 add_339_U1_9 ( .A(xi2_i[56]), .B(xi6_i[56]), .CI(add_339_carry[9]), 
        .CO(add_339_carry[10]), .S(s1_2_i[9]) );
  FA1D0 add_339_U1_8 ( .A(xi2_i[55]), .B(xi6_i[55]), .CI(add_339_carry[8]), 
        .CO(add_339_carry[9]), .S(s1_2_i[8]) );
  FA1D0 add_339_U1_7 ( .A(xi2_i[54]), .B(xi6_i[54]), .CI(add_339_carry[7]), 
        .CO(add_339_carry[8]), .S(s1_2_i[7]) );
  FA1D0 add_339_U1_6 ( .A(xi2_i[53]), .B(xi6_i[53]), .CI(add_339_carry[6]), 
        .CO(add_339_carry[7]), .S(s1_2_i[6]) );
  FA1D0 add_339_U1_5 ( .A(xi2_i[52]), .B(xi6_i[52]), .CI(add_339_carry[5]), 
        .CO(add_339_carry[6]), .S(s1_2_i[5]) );
  FA1D0 add_339_U1_4 ( .A(xi2_i[51]), .B(xi6_i[51]), .CI(add_339_carry[4]), 
        .CO(add_339_carry[5]), .S(s1_2_i[4]) );
  FA1D0 add_339_U1_3 ( .A(xi2_i[50]), .B(xi6_i[50]), .CI(add_339_carry[3]), 
        .CO(add_339_carry[4]), .S(s1_2_i[3]) );
  FA1D0 add_339_U1_2 ( .A(xi2_i[49]), .B(xi6_i[49]), .CI(add_339_carry[2]), 
        .CO(add_339_carry[3]), .S(s1_2_i[2]) );
  FA1D0 add_339_U1_1 ( .A(xi2_i[48]), .B(xi6_i[48]), .CI(add_339_carry[1]), 
        .CO(add_339_carry[2]), .S(s1_2_i[1]) );
  FA1D0 add_331_U1_15 ( .A(xi3_r[62]), .B(xi7_r[62]), .CI(add_331_carry[15]), 
        .CO(add_331_carry[16]), .S(s1_3_r[15]) );
  FA1D0 add_331_U1_14 ( .A(xi3_r[61]), .B(xi7_r[61]), .CI(add_331_carry[14]), 
        .CO(add_331_carry[15]), .S(s1_3_r[14]) );
  FA1D0 add_331_U1_13 ( .A(xi3_r[60]), .B(xi7_r[60]), .CI(add_331_carry[13]), 
        .CO(add_331_carry[14]), .S(s1_3_r[13]) );
  FA1D0 add_331_U1_12 ( .A(xi3_r[59]), .B(xi7_r[59]), .CI(add_331_carry[12]), 
        .CO(add_331_carry[13]), .S(s1_3_r[12]) );
  FA1D0 add_331_U1_11 ( .A(xi3_r[58]), .B(xi7_r[58]), .CI(add_331_carry[11]), 
        .CO(add_331_carry[12]), .S(s1_3_r[11]) );
  FA1D0 add_331_U1_10 ( .A(xi3_r[57]), .B(xi7_r[57]), .CI(add_331_carry[10]), 
        .CO(add_331_carry[11]), .S(s1_3_r[10]) );
  FA1D0 add_331_U1_9 ( .A(xi3_r[56]), .B(xi7_r[56]), .CI(add_331_carry[9]), 
        .CO(add_331_carry[10]), .S(s1_3_r[9]) );
  FA1D0 add_331_U1_8 ( .A(xi3_r[55]), .B(xi7_r[55]), .CI(add_331_carry[8]), 
        .CO(add_331_carry[9]), .S(s1_3_r[8]) );
  FA1D0 add_331_U1_7 ( .A(xi3_r[54]), .B(xi7_r[54]), .CI(add_331_carry[7]), 
        .CO(add_331_carry[8]), .S(s1_3_r[7]) );
  FA1D0 add_331_U1_6 ( .A(xi3_r[53]), .B(xi7_r[53]), .CI(add_331_carry[6]), 
        .CO(add_331_carry[7]), .S(s1_3_r[6]) );
  FA1D0 add_331_U1_5 ( .A(xi3_r[52]), .B(xi7_r[52]), .CI(add_331_carry[5]), 
        .CO(add_331_carry[6]), .S(s1_3_r[5]) );
  FA1D0 add_331_U1_4 ( .A(xi3_r[51]), .B(xi7_r[51]), .CI(add_331_carry[4]), 
        .CO(add_331_carry[5]), .S(s1_3_r[4]) );
  FA1D0 add_331_U1_3 ( .A(xi3_r[50]), .B(xi7_r[50]), .CI(add_331_carry[3]), 
        .CO(add_331_carry[4]), .S(s1_3_r[3]) );
  FA1D0 add_331_U1_2 ( .A(xi3_r[49]), .B(xi7_r[49]), .CI(add_331_carry[2]), 
        .CO(add_331_carry[3]), .S(s1_3_r[2]) );
  FA1D0 add_331_U1_1 ( .A(xi3_r[48]), .B(xi7_r[48]), .CI(add_331_carry[1]), 
        .CO(add_331_carry[2]), .S(s1_3_r[1]) );
  FA1D0 add_340_U1_15 ( .A(xi3_i[62]), .B(xi7_i[62]), .CI(add_340_carry[15]), 
        .CO(add_340_carry[16]), .S(s1_3_i[15]) );
  FA1D0 add_340_U1_14 ( .A(xi3_i[61]), .B(xi7_i[61]), .CI(add_340_carry[14]), 
        .CO(add_340_carry[15]), .S(s1_3_i[14]) );
  FA1D0 add_340_U1_13 ( .A(xi3_i[60]), .B(xi7_i[60]), .CI(add_340_carry[13]), 
        .CO(add_340_carry[14]), .S(s1_3_i[13]) );
  FA1D0 add_340_U1_12 ( .A(xi3_i[59]), .B(xi7_i[59]), .CI(add_340_carry[12]), 
        .CO(add_340_carry[13]), .S(s1_3_i[12]) );
  FA1D0 add_340_U1_11 ( .A(xi3_i[58]), .B(xi7_i[58]), .CI(add_340_carry[11]), 
        .CO(add_340_carry[12]), .S(s1_3_i[11]) );
  FA1D0 add_340_U1_10 ( .A(xi3_i[57]), .B(xi7_i[57]), .CI(add_340_carry[10]), 
        .CO(add_340_carry[11]), .S(s1_3_i[10]) );
  FA1D0 add_340_U1_9 ( .A(xi3_i[56]), .B(xi7_i[56]), .CI(add_340_carry[9]), 
        .CO(add_340_carry[10]), .S(s1_3_i[9]) );
  FA1D0 add_340_U1_8 ( .A(xi3_i[55]), .B(xi7_i[55]), .CI(add_340_carry[8]), 
        .CO(add_340_carry[9]), .S(s1_3_i[8]) );
  FA1D0 add_340_U1_7 ( .A(xi3_i[54]), .B(xi7_i[54]), .CI(add_340_carry[7]), 
        .CO(add_340_carry[8]), .S(s1_3_i[7]) );
  FA1D0 add_340_U1_6 ( .A(xi3_i[53]), .B(xi7_i[53]), .CI(add_340_carry[6]), 
        .CO(add_340_carry[7]), .S(s1_3_i[6]) );
  FA1D0 add_340_U1_5 ( .A(xi3_i[52]), .B(xi7_i[52]), .CI(add_340_carry[5]), 
        .CO(add_340_carry[6]), .S(s1_3_i[5]) );
  FA1D0 add_340_U1_4 ( .A(xi3_i[51]), .B(xi7_i[51]), .CI(add_340_carry[4]), 
        .CO(add_340_carry[5]), .S(s1_3_i[4]) );
  FA1D0 add_340_U1_3 ( .A(xi3_i[50]), .B(xi7_i[50]), .CI(add_340_carry[3]), 
        .CO(add_340_carry[4]), .S(s1_3_i[3]) );
  FA1D0 add_340_U1_2 ( .A(xi3_i[49]), .B(xi7_i[49]), .CI(add_340_carry[2]), 
        .CO(add_340_carry[3]), .S(s1_3_i[2]) );
  FA1D0 add_340_U1_1 ( .A(xi3_i[48]), .B(xi7_i[48]), .CI(add_340_carry[1]), 
        .CO(add_340_carry[2]), .S(s1_3_i[1]) );
  FA1D0 sub_332_U2_15 ( .A(xi0_r[62]), .B(n1177), .CI(sub_332_carry[15]), .CO(
        sub_332_carry[16]), .S(s1_4_r[15]) );
  FA1D0 sub_332_U2_14 ( .A(xi0_r[61]), .B(n1178), .CI(sub_332_carry[14]), .CO(
        sub_332_carry[15]), .S(s1_4_r[14]) );
  FA1D0 sub_332_U2_13 ( .A(xi0_r[60]), .B(n1179), .CI(sub_332_carry[13]), .CO(
        sub_332_carry[14]), .S(s1_4_r[13]) );
  FA1D0 sub_332_U2_12 ( .A(xi0_r[59]), .B(n1180), .CI(sub_332_carry[12]), .CO(
        sub_332_carry[13]), .S(s1_4_r[12]) );
  FA1D0 sub_332_U2_11 ( .A(xi0_r[58]), .B(n1181), .CI(sub_332_carry[11]), .CO(
        sub_332_carry[12]), .S(s1_4_r[11]) );
  FA1D0 sub_332_U2_10 ( .A(xi0_r[57]), .B(n1182), .CI(sub_332_carry[10]), .CO(
        sub_332_carry[11]), .S(s1_4_r[10]) );
  FA1D0 sub_332_U2_9 ( .A(xi0_r[56]), .B(n1183), .CI(sub_332_carry[9]), .CO(
        sub_332_carry[10]), .S(s1_4_r[9]) );
  FA1D0 sub_332_U2_8 ( .A(xi0_r[55]), .B(n1184), .CI(sub_332_carry[8]), .CO(
        sub_332_carry[9]), .S(s1_4_r[8]) );
  FA1D0 sub_332_U2_7 ( .A(xi0_r[54]), .B(n1185), .CI(sub_332_carry[7]), .CO(
        sub_332_carry[8]), .S(s1_4_r[7]) );
  FA1D0 sub_332_U2_6 ( .A(xi0_r[53]), .B(n1186), .CI(sub_332_carry[6]), .CO(
        sub_332_carry[7]), .S(s1_4_r[6]) );
  FA1D0 sub_332_U2_5 ( .A(xi0_r[52]), .B(n1187), .CI(sub_332_carry[5]), .CO(
        sub_332_carry[6]), .S(s1_4_r[5]) );
  FA1D0 sub_332_U2_4 ( .A(xi0_r[51]), .B(n1188), .CI(sub_332_carry[4]), .CO(
        sub_332_carry[5]), .S(s1_4_r[4]) );
  FA1D0 sub_332_U2_3 ( .A(xi0_r[50]), .B(n1189), .CI(sub_332_carry[3]), .CO(
        sub_332_carry[4]), .S(s1_4_r[3]) );
  FA1D0 sub_332_U2_2 ( .A(xi0_r[49]), .B(n1190), .CI(sub_332_carry[2]), .CO(
        sub_332_carry[3]), .S(s1_4_r[2]) );
  FA1D0 sub_332_U2_1 ( .A(xi0_r[48]), .B(n1191), .CI(sub_332_carry[1]), .CO(
        sub_332_carry[2]), .S(s1_4_r[1]) );
  FA1D0 sub_341_U2_15 ( .A(xi0_i[62]), .B(n1307), .CI(sub_341_carry[15]), .CO(
        sub_341_carry[16]), .S(s1_4_i[15]) );
  FA1D0 sub_341_U2_14 ( .A(xi0_i[61]), .B(n1308), .CI(sub_341_carry[14]), .CO(
        sub_341_carry[15]), .S(s1_4_i[14]) );
  FA1D0 sub_341_U2_13 ( .A(xi0_i[60]), .B(n1309), .CI(sub_341_carry[13]), .CO(
        sub_341_carry[14]), .S(s1_4_i[13]) );
  FA1D0 sub_341_U2_12 ( .A(xi0_i[59]), .B(n1310), .CI(sub_341_carry[12]), .CO(
        sub_341_carry[13]), .S(s1_4_i[12]) );
  FA1D0 sub_341_U2_11 ( .A(xi0_i[58]), .B(n1311), .CI(sub_341_carry[11]), .CO(
        sub_341_carry[12]), .S(s1_4_i[11]) );
  FA1D0 sub_341_U2_10 ( .A(xi0_i[57]), .B(n1312), .CI(sub_341_carry[10]), .CO(
        sub_341_carry[11]), .S(s1_4_i[10]) );
  FA1D0 sub_341_U2_9 ( .A(xi0_i[56]), .B(n1313), .CI(sub_341_carry[9]), .CO(
        sub_341_carry[10]), .S(s1_4_i[9]) );
  FA1D0 sub_341_U2_8 ( .A(xi0_i[55]), .B(n1314), .CI(sub_341_carry[8]), .CO(
        sub_341_carry[9]), .S(s1_4_i[8]) );
  FA1D0 sub_341_U2_7 ( .A(xi0_i[54]), .B(n1315), .CI(sub_341_carry[7]), .CO(
        sub_341_carry[8]), .S(s1_4_i[7]) );
  FA1D0 sub_341_U2_6 ( .A(xi0_i[53]), .B(n1316), .CI(sub_341_carry[6]), .CO(
        sub_341_carry[7]), .S(s1_4_i[6]) );
  FA1D0 sub_341_U2_5 ( .A(xi0_i[52]), .B(n1317), .CI(sub_341_carry[5]), .CO(
        sub_341_carry[6]), .S(s1_4_i[5]) );
  FA1D0 sub_341_U2_4 ( .A(xi0_i[51]), .B(n1318), .CI(sub_341_carry[4]), .CO(
        sub_341_carry[5]), .S(s1_4_i[4]) );
  FA1D0 sub_341_U2_3 ( .A(xi0_i[50]), .B(n1319), .CI(sub_341_carry[3]), .CO(
        sub_341_carry[4]), .S(s1_4_i[3]) );
  FA1D0 sub_341_U2_2 ( .A(xi0_i[49]), .B(n1320), .CI(sub_341_carry[2]), .CO(
        sub_341_carry[3]), .S(s1_4_i[2]) );
  FA1D0 sub_341_U2_1 ( .A(xi0_i[48]), .B(n1321), .CI(sub_341_carry[1]), .CO(
        sub_341_carry[2]), .S(s1_4_i[1]) );
  FA1D0 sub_343_U2_15 ( .A(xi2_i[62]), .B(n1339), .CI(sub_343_carry[15]), .CO(
        sub_343_carry[16]), .S(s1_6_i[15]) );
  FA1D0 sub_343_U2_14 ( .A(xi2_i[61]), .B(n1340), .CI(sub_343_carry[14]), .CO(
        sub_343_carry[15]), .S(s1_6_i[14]) );
  FA1D0 sub_343_U2_13 ( .A(xi2_i[60]), .B(n1341), .CI(sub_343_carry[13]), .CO(
        sub_343_carry[14]), .S(s1_6_i[13]) );
  FA1D0 sub_343_U2_12 ( .A(xi2_i[59]), .B(n1342), .CI(sub_343_carry[12]), .CO(
        sub_343_carry[13]), .S(s1_6_i[12]) );
  FA1D0 sub_343_U2_11 ( .A(xi2_i[58]), .B(n1343), .CI(sub_343_carry[11]), .CO(
        sub_343_carry[12]), .S(s1_6_i[11]) );
  FA1D0 sub_343_U2_10 ( .A(xi2_i[57]), .B(n1344), .CI(sub_343_carry[10]), .CO(
        sub_343_carry[11]), .S(s1_6_i[10]) );
  FA1D0 sub_343_U2_9 ( .A(xi2_i[56]), .B(n1345), .CI(sub_343_carry[9]), .CO(
        sub_343_carry[10]), .S(s1_6_i[9]) );
  FA1D0 sub_343_U2_8 ( .A(xi2_i[55]), .B(n1346), .CI(sub_343_carry[8]), .CO(
        sub_343_carry[9]), .S(s1_6_i[8]) );
  FA1D0 sub_343_U2_7 ( .A(xi2_i[54]), .B(n1347), .CI(sub_343_carry[7]), .CO(
        sub_343_carry[8]), .S(s1_6_i[7]) );
  FA1D0 sub_343_U2_6 ( .A(xi2_i[53]), .B(n1348), .CI(sub_343_carry[6]), .CO(
        sub_343_carry[7]), .S(s1_6_i[6]) );
  FA1D0 sub_343_U2_5 ( .A(xi2_i[52]), .B(n1349), .CI(sub_343_carry[5]), .CO(
        sub_343_carry[6]), .S(s1_6_i[5]) );
  FA1D0 sub_343_U2_4 ( .A(xi2_i[51]), .B(n1350), .CI(sub_343_carry[4]), .CO(
        sub_343_carry[5]), .S(s1_6_i[4]) );
  FA1D0 sub_343_U2_3 ( .A(xi2_i[50]), .B(n1351), .CI(sub_343_carry[3]), .CO(
        sub_343_carry[4]), .S(s1_6_i[3]) );
  FA1D0 sub_343_U2_2 ( .A(xi2_i[49]), .B(n1352), .CI(sub_343_carry[2]), .CO(
        sub_343_carry[3]), .S(s1_6_i[2]) );
  FA1D0 sub_343_U2_1 ( .A(xi2_i[48]), .B(n1353), .CI(sub_343_carry[1]), .CO(
        sub_343_carry[2]), .S(s1_6_i[1]) );
  FA1D0 sub_334_U2_1 ( .A(xi2_r[48]), .B(n1223), .CI(sub_334_carry[1]), .CO(
        sub_334_carry[2]), .S(s1_6_tmp_i[0]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_1 ( .A(xo7_r_w_d1r[1]), .B(n1602), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[1]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[2]), .S(dp_cluster_4_s2_7_r[9])
         );
  FA1D0 sub_365_U2_1 ( .A(xo5_i_w_d1r[1]), .B(n1684), .CI(sub_365_carry[1]), 
        .CO(sub_365_carry[2]), .S(s2_7_i[1]) );
  FA1D0 add_350_U1_1 ( .A(xo1_r_w_d1r[1]), .B(xo3_r_w_d1r[1]), .CI(n922), .CO(
        add_350_carry[2]), .S(s2_1_r[1]) );
  FA1D0 add_359_U1_1 ( .A(xo1_i_w_d1r[1]), .B(xo3_i_w_d1r[1]), .CI(n920), .CO(
        add_359_carry[2]), .S(s2_1_i[1]) );
  FA1D0 sub_361_U2_1 ( .A(xo1_i_w_d1r[1]), .B(n1556), .CI(sub_361_carry[1]), 
        .CO(sub_361_carry[2]), .S(s2_3_i[1]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_1 ( .A(xo3_r_w_d1r[1]), .B(n1474), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[1]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[2]), .S(dp_cluster_5_s2_3_r[9])
         );
  FA1D0 add_354_U1_1 ( .A(xo5_r_w_d1r[1]), .B(xo7_r_w_d1r[1]), .CI(n921), .CO(
        add_354_carry[2]), .S(s2_5_r[1]) );
  FA1D0 add_363_U1_1 ( .A(xo5_i_w_d1r[1]), .B(xo7_i_w_d1r[1]), .CI(n919), .CO(
        add_363_carry[2]), .S(s2_5_i[1]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_13 ( .A(xo7_r_w_d1r[13]), .B(n1566), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[13]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[14]), .S(dp_cluster_4_s2_7_r[12]) );
  FA1D0 sub_364_U2_13 ( .A(xo4_i_w_d1r[13]), .B(n1656), .CI(sub_364_carry[13]), 
        .CO(sub_364_carry[14]), .S(s2_6_i[13]) );
  FA1D0 sub_365_U2_13 ( .A(xo5_i_w_d1r[13]), .B(n1672), .CI(sub_365_carry[13]), 
        .CO(sub_365_carry[14]), .S(s2_7_i[13]) );
  FA1D0 sub_355_U2_13 ( .A(xo4_r_w_d1r[13]), .B(n1640), .CI(sub_355_carry[13]), 
        .CO(sub_355_carry[14]), .S(s2_6_r[13]) );
  FA1D0 add_349_U1_13 ( .A(xo0_r_w_d1r[13]), .B(xo2_r_w_d1r[13]), .CI(
        add_349_carry[13]), .CO(add_349_carry[14]), .S(s2_0_r[13]) );
  FA1D0 add_358_U1_13 ( .A(xo0_i_w_d1r[13]), .B(xo2_i_w_d1r[13]), .CI(
        add_358_carry[13]), .CO(add_358_carry[14]), .S(s2_0_i[13]) );
  FA1D0 sub_351_U2_13 ( .A(xo0_r_w_d1r[13]), .B(n1512), .CI(sub_351_carry[13]), 
        .CO(sub_351_carry[14]), .S(s2_2_r[13]) );
  FA1D0 sub_360_U2_13 ( .A(xo0_i_w_d1r[13]), .B(n1528), .CI(sub_360_carry[13]), 
        .CO(sub_360_carry[14]), .S(s2_2_i[13]) );
  FA1D0 add_353_U1_13 ( .A(xo4_r_w_d1r[13]), .B(xo6_r_w_d1r[13]), .CI(
        add_353_carry[13]), .CO(add_353_carry[14]), .S(s2_4_r[13]) );
  FA1D0 add_362_U1_13 ( .A(xo4_i_w_d1r[13]), .B(xo6_i_w_d1r[13]), .CI(
        add_362_carry[13]), .CO(add_362_carry[14]), .S(s2_4_i[13]) );
  FA1D0 sub_334_U2_15 ( .A(xi2_r[62]), .B(n1209), .CI(sub_334_carry[15]), .CO(
        sub_334_carry[16]), .S(s1_6_r[15]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_12 ( .A(xo7_r_w_d1r[12]), .B(n1569), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[12]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[13]), .S(dp_cluster_4_s2_7_r[13]) );
  FA1D0 sub_364_U2_12 ( .A(xo4_i_w_d1r[12]), .B(n1657), .CI(sub_364_carry[12]), 
        .CO(sub_364_carry[13]), .S(s2_6_i[12]) );
  FA1D0 sub_365_U2_12 ( .A(xo5_i_w_d1r[12]), .B(n1673), .CI(sub_365_carry[12]), 
        .CO(sub_365_carry[13]), .S(s2_7_i[12]) );
  FA1D0 sub_355_U2_12 ( .A(xo4_r_w_d1r[12]), .B(n1641), .CI(sub_355_carry[12]), 
        .CO(sub_355_carry[13]), .S(s2_6_r[12]) );
  FA1D0 add_349_U1_12 ( .A(xo0_r_w_d1r[12]), .B(xo2_r_w_d1r[12]), .CI(
        add_349_carry[12]), .CO(add_349_carry[13]), .S(s2_0_r[12]) );
  FA1D0 add_358_U1_12 ( .A(xo0_i_w_d1r[12]), .B(xo2_i_w_d1r[12]), .CI(
        add_358_carry[12]), .CO(add_358_carry[13]), .S(s2_0_i[12]) );
  FA1D0 add_350_U1_13 ( .A(xo1_r_w_d1r[13]), .B(xo3_r_w_d1r[13]), .CI(
        add_350_carry[13]), .CO(add_350_carry[14]), .S(s2_1_r[13]) );
  FA1D0 add_359_U1_13 ( .A(xo1_i_w_d1r[13]), .B(xo3_i_w_d1r[13]), .CI(
        add_359_carry[13]), .CO(add_359_carry[14]), .S(s2_1_i[13]) );
  FA1D0 sub_351_U2_12 ( .A(xo0_r_w_d1r[12]), .B(n1513), .CI(sub_351_carry[12]), 
        .CO(sub_351_carry[13]), .S(s2_2_r[12]) );
  FA1D0 sub_360_U2_12 ( .A(xo0_i_w_d1r[12]), .B(n1529), .CI(sub_360_carry[12]), 
        .CO(sub_360_carry[13]), .S(s2_2_i[12]) );
  FA1D0 sub_361_U2_13 ( .A(xo1_i_w_d1r[13]), .B(n1544), .CI(sub_361_carry[13]), 
        .CO(sub_361_carry[14]), .S(s2_3_i[13]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_13 ( .A(xo3_r_w_d1r[13]), .B(n1438), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[13]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[14]), .S(dp_cluster_5_s2_3_r[12]) );
  FA1D0 add_353_U1_12 ( .A(xo4_r_w_d1r[12]), .B(xo6_r_w_d1r[12]), .CI(
        add_353_carry[12]), .CO(add_353_carry[13]), .S(s2_4_r[12]) );
  FA1D0 add_362_U1_12 ( .A(xo4_i_w_d1r[12]), .B(xo6_i_w_d1r[12]), .CI(
        add_362_carry[12]), .CO(add_362_carry[13]), .S(s2_4_i[12]) );
  FA1D0 add_354_U1_13 ( .A(xo5_r_w_d1r[13]), .B(xo7_r_w_d1r[13]), .CI(
        add_354_carry[13]), .CO(add_354_carry[14]), .S(s2_5_r[13]) );
  FA1D0 add_363_U1_13 ( .A(xo5_i_w_d1r[13]), .B(xo7_i_w_d1r[13]), .CI(
        add_363_carry[13]), .CO(add_363_carry[14]), .S(s2_5_i[13]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_11 ( .A(xo7_r_w_d1r[11]), .B(n1572), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[11]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[12]), .S(dp_cluster_4_s2_7_r[14]) );
  FA1D0 sub_364_U2_11 ( .A(xo4_i_w_d1r[11]), .B(n1658), .CI(sub_364_carry[11]), 
        .CO(sub_364_carry[12]), .S(s2_6_i[11]) );
  FA1D0 sub_365_U2_11 ( .A(xo5_i_w_d1r[11]), .B(n1674), .CI(sub_365_carry[11]), 
        .CO(sub_365_carry[12]), .S(s2_7_i[11]) );
  FA1D0 sub_355_U2_11 ( .A(xo4_r_w_d1r[11]), .B(n1642), .CI(sub_355_carry[11]), 
        .CO(sub_355_carry[12]), .S(s2_6_r[11]) );
  FA1D0 add_349_U1_11 ( .A(xo0_r_w_d1r[11]), .B(xo2_r_w_d1r[11]), .CI(
        add_349_carry[11]), .CO(add_349_carry[12]), .S(s2_0_r[11]) );
  FA1D0 add_358_U1_11 ( .A(xo0_i_w_d1r[11]), .B(xo2_i_w_d1r[11]), .CI(
        add_358_carry[11]), .CO(add_358_carry[12]), .S(s2_0_i[11]) );
  FA1D0 add_350_U1_12 ( .A(xo1_r_w_d1r[12]), .B(xo3_r_w_d1r[12]), .CI(
        add_350_carry[12]), .CO(add_350_carry[13]), .S(s2_1_r[12]) );
  FA1D0 add_359_U1_12 ( .A(xo1_i_w_d1r[12]), .B(xo3_i_w_d1r[12]), .CI(
        add_359_carry[12]), .CO(add_359_carry[13]), .S(s2_1_i[12]) );
  FA1D0 sub_351_U2_11 ( .A(xo0_r_w_d1r[11]), .B(n1514), .CI(sub_351_carry[11]), 
        .CO(sub_351_carry[12]), .S(s2_2_r[11]) );
  FA1D0 sub_360_U2_11 ( .A(xo0_i_w_d1r[11]), .B(n1530), .CI(sub_360_carry[11]), 
        .CO(sub_360_carry[12]), .S(s2_2_i[11]) );
  FA1D0 sub_361_U2_12 ( .A(xo1_i_w_d1r[12]), .B(n1545), .CI(sub_361_carry[12]), 
        .CO(sub_361_carry[13]), .S(s2_3_i[12]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_12 ( .A(xo3_r_w_d1r[12]), .B(n1441), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[12]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[13]), .S(dp_cluster_5_s2_3_r[13]) );
  FA1D0 add_353_U1_11 ( .A(xo4_r_w_d1r[11]), .B(xo6_r_w_d1r[11]), .CI(
        add_353_carry[11]), .CO(add_353_carry[12]), .S(s2_4_r[11]) );
  FA1D0 add_362_U1_11 ( .A(xo4_i_w_d1r[11]), .B(xo6_i_w_d1r[11]), .CI(
        add_362_carry[11]), .CO(add_362_carry[12]), .S(s2_4_i[11]) );
  FA1D0 add_354_U1_12 ( .A(xo5_r_w_d1r[12]), .B(xo7_r_w_d1r[12]), .CI(
        add_354_carry[12]), .CO(add_354_carry[13]), .S(s2_5_r[12]) );
  FA1D0 add_363_U1_12 ( .A(xo5_i_w_d1r[12]), .B(xo7_i_w_d1r[12]), .CI(
        add_363_carry[12]), .CO(add_363_carry[13]), .S(s2_5_i[12]) );
  FA1D0 sub_334_U2_14 ( .A(xi2_r[61]), .B(n1210), .CI(sub_334_carry[14]), .CO(
        sub_334_carry[15]), .S(s1_6_r[14]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_10 ( .A(xo7_r_w_d1r[10]), .B(n1575), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[10]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[11]), .S(dp_cluster_4_s2_7_r[15]) );
  FA1D0 sub_364_U2_10 ( .A(xo4_i_w_d1r[10]), .B(n1659), .CI(sub_364_carry[10]), 
        .CO(sub_364_carry[11]), .S(s2_6_i[10]) );
  FA1D0 sub_365_U2_10 ( .A(xo5_i_w_d1r[10]), .B(n1675), .CI(sub_365_carry[10]), 
        .CO(sub_365_carry[11]), .S(s2_7_i[10]) );
  FA1D0 sub_355_U2_10 ( .A(xo4_r_w_d1r[10]), .B(n1643), .CI(sub_355_carry[10]), 
        .CO(sub_355_carry[11]), .S(s2_6_r[10]) );
  FA1D0 add_349_U1_10 ( .A(xo0_r_w_d1r[10]), .B(xo2_r_w_d1r[10]), .CI(
        add_349_carry[10]), .CO(add_349_carry[11]), .S(s2_0_r[10]) );
  FA1D0 add_358_U1_10 ( .A(xo0_i_w_d1r[10]), .B(xo2_i_w_d1r[10]), .CI(
        add_358_carry[10]), .CO(add_358_carry[11]), .S(s2_0_i[10]) );
  FA1D0 add_350_U1_11 ( .A(xo1_r_w_d1r[11]), .B(xo3_r_w_d1r[11]), .CI(
        add_350_carry[11]), .CO(add_350_carry[12]), .S(s2_1_r[11]) );
  FA1D0 add_359_U1_11 ( .A(xo1_i_w_d1r[11]), .B(xo3_i_w_d1r[11]), .CI(
        add_359_carry[11]), .CO(add_359_carry[12]), .S(s2_1_i[11]) );
  FA1D0 sub_351_U2_10 ( .A(xo0_r_w_d1r[10]), .B(n1515), .CI(sub_351_carry[10]), 
        .CO(sub_351_carry[11]), .S(s2_2_r[10]) );
  FA1D0 sub_360_U2_10 ( .A(xo0_i_w_d1r[10]), .B(n1531), .CI(sub_360_carry[10]), 
        .CO(sub_360_carry[11]), .S(s2_2_i[10]) );
  FA1D0 sub_361_U2_11 ( .A(xo1_i_w_d1r[11]), .B(n1546), .CI(sub_361_carry[11]), 
        .CO(sub_361_carry[12]), .S(s2_3_i[11]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_11 ( .A(xo3_r_w_d1r[11]), .B(n1444), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[11]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[12]), .S(dp_cluster_5_s2_3_r[14]) );
  FA1D0 add_353_U1_10 ( .A(xo4_r_w_d1r[10]), .B(xo6_r_w_d1r[10]), .CI(
        add_353_carry[10]), .CO(add_353_carry[11]), .S(s2_4_r[10]) );
  FA1D0 add_362_U1_10 ( .A(xo4_i_w_d1r[10]), .B(xo6_i_w_d1r[10]), .CI(
        add_362_carry[10]), .CO(add_362_carry[11]), .S(s2_4_i[10]) );
  FA1D0 add_354_U1_11 ( .A(xo5_r_w_d1r[11]), .B(xo7_r_w_d1r[11]), .CI(
        add_354_carry[11]), .CO(add_354_carry[12]), .S(s2_5_r[11]) );
  FA1D0 add_363_U1_11 ( .A(xo5_i_w_d1r[11]), .B(xo7_i_w_d1r[11]), .CI(
        add_363_carry[11]), .CO(add_363_carry[12]), .S(s2_5_i[11]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_9 ( .A(xo7_r_w_d1r[9]), .B(n1578), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[9]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[10]), .S(dp_cluster_4_s2_7_r[1])
         );
  FA1D0 sub_364_U2_9 ( .A(xo4_i_w_d1r[9]), .B(n1660), .CI(sub_364_carry[9]), 
        .CO(sub_364_carry[10]), .S(s2_6_i[9]) );
  FA1D0 sub_365_U2_9 ( .A(xo5_i_w_d1r[9]), .B(n1676), .CI(sub_365_carry[9]), 
        .CO(sub_365_carry[10]), .S(s2_7_i[9]) );
  FA1D0 sub_355_U2_9 ( .A(xo4_r_w_d1r[9]), .B(n1644), .CI(sub_355_carry[9]), 
        .CO(sub_355_carry[10]), .S(s2_6_r[9]) );
  FA1D0 add_349_U1_9 ( .A(xo0_r_w_d1r[9]), .B(xo2_r_w_d1r[9]), .CI(
        add_349_carry[9]), .CO(add_349_carry[10]), .S(s2_0_r[9]) );
  FA1D0 add_358_U1_9 ( .A(xo0_i_w_d1r[9]), .B(xo2_i_w_d1r[9]), .CI(
        add_358_carry[9]), .CO(add_358_carry[10]), .S(s2_0_i[9]) );
  FA1D0 add_350_U1_10 ( .A(xo1_r_w_d1r[10]), .B(xo3_r_w_d1r[10]), .CI(
        add_350_carry[10]), .CO(add_350_carry[11]), .S(s2_1_r[10]) );
  FA1D0 add_359_U1_10 ( .A(xo1_i_w_d1r[10]), .B(xo3_i_w_d1r[10]), .CI(
        add_359_carry[10]), .CO(add_359_carry[11]), .S(s2_1_i[10]) );
  FA1D0 sub_351_U2_9 ( .A(xo0_r_w_d1r[9]), .B(n1516), .CI(sub_351_carry[9]), 
        .CO(sub_351_carry[10]), .S(s2_2_r[9]) );
  FA1D0 sub_360_U2_9 ( .A(xo0_i_w_d1r[9]), .B(n1532), .CI(sub_360_carry[9]), 
        .CO(sub_360_carry[10]), .S(s2_2_i[9]) );
  FA1D0 sub_361_U2_10 ( .A(xo1_i_w_d1r[10]), .B(n1547), .CI(sub_361_carry[10]), 
        .CO(sub_361_carry[11]), .S(s2_3_i[10]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_10 ( .A(xo3_r_w_d1r[10]), .B(n1447), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[10]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[11]), .S(dp_cluster_5_s2_3_r[15]) );
  FA1D0 add_353_U1_9 ( .A(xo4_r_w_d1r[9]), .B(xo6_r_w_d1r[9]), .CI(
        add_353_carry[9]), .CO(add_353_carry[10]), .S(s2_4_r[9]) );
  FA1D0 add_362_U1_9 ( .A(xo4_i_w_d1r[9]), .B(xo6_i_w_d1r[9]), .CI(
        add_362_carry[9]), .CO(add_362_carry[10]), .S(s2_4_i[9]) );
  FA1D0 add_354_U1_10 ( .A(xo5_r_w_d1r[10]), .B(xo7_r_w_d1r[10]), .CI(
        add_354_carry[10]), .CO(add_354_carry[11]), .S(s2_5_r[10]) );
  FA1D0 add_363_U1_10 ( .A(xo5_i_w_d1r[10]), .B(xo7_i_w_d1r[10]), .CI(
        add_363_carry[10]), .CO(add_363_carry[11]), .S(s2_5_i[10]) );
  FA1D0 sub_334_U2_13 ( .A(xi2_r[60]), .B(n1211), .CI(sub_334_carry[13]), .CO(
        sub_334_carry[14]), .S(s1_6_r[13]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_8 ( .A(xo7_r_w_d1r[8]), .B(n1581), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[8]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[9]), .S(dp_cluster_4_s2_7_r[2])
         );
  FA1D0 sub_364_U2_8 ( .A(xo4_i_w_d1r[8]), .B(n1661), .CI(sub_364_carry[8]), 
        .CO(sub_364_carry[9]), .S(s2_6_i[8]) );
  FA1D0 sub_365_U2_8 ( .A(xo5_i_w_d1r[8]), .B(n1677), .CI(sub_365_carry[8]), 
        .CO(sub_365_carry[9]), .S(s2_7_i[8]) );
  FA1D0 sub_355_U2_8 ( .A(xo4_r_w_d1r[8]), .B(n1645), .CI(sub_355_carry[8]), 
        .CO(sub_355_carry[9]), .S(s2_6_r[8]) );
  FA1D0 add_349_U1_8 ( .A(xo0_r_w_d1r[8]), .B(xo2_r_w_d1r[8]), .CI(
        add_349_carry[8]), .CO(add_349_carry[9]), .S(s2_0_r[8]) );
  FA1D0 add_358_U1_8 ( .A(xo0_i_w_d1r[8]), .B(xo2_i_w_d1r[8]), .CI(
        add_358_carry[8]), .CO(add_358_carry[9]), .S(s2_0_i[8]) );
  FA1D0 add_350_U1_9 ( .A(xo1_r_w_d1r[9]), .B(xo3_r_w_d1r[9]), .CI(
        add_350_carry[9]), .CO(add_350_carry[10]), .S(s2_1_r[9]) );
  FA1D0 add_359_U1_9 ( .A(xo1_i_w_d1r[9]), .B(xo3_i_w_d1r[9]), .CI(
        add_359_carry[9]), .CO(add_359_carry[10]), .S(s2_1_i[9]) );
  FA1D0 sub_351_U2_8 ( .A(xo0_r_w_d1r[8]), .B(n1517), .CI(sub_351_carry[8]), 
        .CO(sub_351_carry[9]), .S(s2_2_r[8]) );
  FA1D0 sub_360_U2_8 ( .A(xo0_i_w_d1r[8]), .B(n1533), .CI(sub_360_carry[8]), 
        .CO(sub_360_carry[9]), .S(s2_2_i[8]) );
  FA1D0 sub_361_U2_9 ( .A(xo1_i_w_d1r[9]), .B(n1548), .CI(sub_361_carry[9]), 
        .CO(sub_361_carry[10]), .S(s2_3_i[9]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_9 ( .A(xo3_r_w_d1r[9]), .B(n1450), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[9]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[10]), .S(dp_cluster_5_s2_3_r[1])
         );
  FA1D0 add_353_U1_8 ( .A(xo4_r_w_d1r[8]), .B(xo6_r_w_d1r[8]), .CI(
        add_353_carry[8]), .CO(add_353_carry[9]), .S(s2_4_r[8]) );
  FA1D0 add_362_U1_8 ( .A(xo4_i_w_d1r[8]), .B(xo6_i_w_d1r[8]), .CI(
        add_362_carry[8]), .CO(add_362_carry[9]), .S(s2_4_i[8]) );
  FA1D0 add_354_U1_9 ( .A(xo5_r_w_d1r[9]), .B(xo7_r_w_d1r[9]), .CI(
        add_354_carry[9]), .CO(add_354_carry[10]), .S(s2_5_r[9]) );
  FA1D0 add_363_U1_9 ( .A(xo5_i_w_d1r[9]), .B(xo7_i_w_d1r[9]), .CI(
        add_363_carry[9]), .CO(add_363_carry[10]), .S(s2_5_i[9]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_7 ( .A(xo7_r_w_d1r[7]), .B(n1584), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[7]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[8]), .S(dp_cluster_4_s2_7_r[3])
         );
  FA1D0 sub_364_U2_7 ( .A(xo4_i_w_d1r[7]), .B(n1662), .CI(sub_364_carry[7]), 
        .CO(sub_364_carry[8]), .S(s2_6_i[7]) );
  FA1D0 sub_365_U2_7 ( .A(xo5_i_w_d1r[7]), .B(n1678), .CI(sub_365_carry[7]), 
        .CO(sub_365_carry[8]), .S(s2_7_i[7]) );
  FA1D0 sub_355_U2_7 ( .A(xo4_r_w_d1r[7]), .B(n1646), .CI(sub_355_carry[7]), 
        .CO(sub_355_carry[8]), .S(s2_6_r[7]) );
  FA1D0 add_349_U1_7 ( .A(xo0_r_w_d1r[7]), .B(xo2_r_w_d1r[7]), .CI(
        add_349_carry[7]), .CO(add_349_carry[8]), .S(s2_0_r[7]) );
  FA1D0 add_358_U1_7 ( .A(xo0_i_w_d1r[7]), .B(xo2_i_w_d1r[7]), .CI(
        add_358_carry[7]), .CO(add_358_carry[8]), .S(s2_0_i[7]) );
  FA1D0 add_350_U1_8 ( .A(xo1_r_w_d1r[8]), .B(xo3_r_w_d1r[8]), .CI(
        add_350_carry[8]), .CO(add_350_carry[9]), .S(s2_1_r[8]) );
  FA1D0 add_359_U1_8 ( .A(xo1_i_w_d1r[8]), .B(xo3_i_w_d1r[8]), .CI(
        add_359_carry[8]), .CO(add_359_carry[9]), .S(s2_1_i[8]) );
  FA1D0 sub_351_U2_7 ( .A(xo0_r_w_d1r[7]), .B(n1518), .CI(sub_351_carry[7]), 
        .CO(sub_351_carry[8]), .S(s2_2_r[7]) );
  FA1D0 sub_360_U2_7 ( .A(xo0_i_w_d1r[7]), .B(n1534), .CI(sub_360_carry[7]), 
        .CO(sub_360_carry[8]), .S(s2_2_i[7]) );
  FA1D0 sub_361_U2_8 ( .A(xo1_i_w_d1r[8]), .B(n1549), .CI(sub_361_carry[8]), 
        .CO(sub_361_carry[9]), .S(s2_3_i[8]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_8 ( .A(xo3_r_w_d1r[8]), .B(n1453), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[8]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[9]), .S(dp_cluster_5_s2_3_r[2])
         );
  FA1D0 add_353_U1_7 ( .A(xo4_r_w_d1r[7]), .B(xo6_r_w_d1r[7]), .CI(
        add_353_carry[7]), .CO(add_353_carry[8]), .S(s2_4_r[7]) );
  FA1D0 add_362_U1_7 ( .A(xo4_i_w_d1r[7]), .B(xo6_i_w_d1r[7]), .CI(
        add_362_carry[7]), .CO(add_362_carry[8]), .S(s2_4_i[7]) );
  FA1D0 add_354_U1_8 ( .A(xo5_r_w_d1r[8]), .B(xo7_r_w_d1r[8]), .CI(
        add_354_carry[8]), .CO(add_354_carry[9]), .S(s2_5_r[8]) );
  FA1D0 add_363_U1_8 ( .A(xo5_i_w_d1r[8]), .B(xo7_i_w_d1r[8]), .CI(
        add_363_carry[8]), .CO(add_363_carry[9]), .S(s2_5_i[8]) );
  FA1D0 sub_334_U2_12 ( .A(xi2_r[59]), .B(n1212), .CI(sub_334_carry[12]), .CO(
        sub_334_carry[13]), .S(s1_6_r[12]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_6 ( .A(xo7_r_w_d1r[6]), .B(n1587), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[6]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[7]), .S(dp_cluster_4_s2_7_r[4])
         );
  FA1D0 sub_364_U2_6 ( .A(xo4_i_w_d1r[6]), .B(n1663), .CI(sub_364_carry[6]), 
        .CO(sub_364_carry[7]), .S(s2_6_i[6]) );
  FA1D0 sub_365_U2_6 ( .A(xo5_i_w_d1r[6]), .B(n1679), .CI(sub_365_carry[6]), 
        .CO(sub_365_carry[7]), .S(s2_7_i[6]) );
  FA1D0 sub_355_U2_6 ( .A(xo4_r_w_d1r[6]), .B(n1647), .CI(sub_355_carry[6]), 
        .CO(sub_355_carry[7]), .S(s2_6_r[6]) );
  FA1D0 add_349_U1_6 ( .A(xo0_r_w_d1r[6]), .B(xo2_r_w_d1r[6]), .CI(
        add_349_carry[6]), .CO(add_349_carry[7]), .S(s2_0_r[6]) );
  FA1D0 add_358_U1_6 ( .A(xo0_i_w_d1r[6]), .B(xo2_i_w_d1r[6]), .CI(
        add_358_carry[6]), .CO(add_358_carry[7]), .S(s2_0_i[6]) );
  FA1D0 add_350_U1_7 ( .A(xo1_r_w_d1r[7]), .B(xo3_r_w_d1r[7]), .CI(
        add_350_carry[7]), .CO(add_350_carry[8]), .S(s2_1_r[7]) );
  FA1D0 add_359_U1_7 ( .A(xo1_i_w_d1r[7]), .B(xo3_i_w_d1r[7]), .CI(
        add_359_carry[7]), .CO(add_359_carry[8]), .S(s2_1_i[7]) );
  FA1D0 sub_351_U2_6 ( .A(xo0_r_w_d1r[6]), .B(n1519), .CI(sub_351_carry[6]), 
        .CO(sub_351_carry[7]), .S(s2_2_r[6]) );
  FA1D0 sub_360_U2_6 ( .A(xo0_i_w_d1r[6]), .B(n1535), .CI(sub_360_carry[6]), 
        .CO(sub_360_carry[7]), .S(s2_2_i[6]) );
  FA1D0 sub_361_U2_7 ( .A(xo1_i_w_d1r[7]), .B(n1550), .CI(sub_361_carry[7]), 
        .CO(sub_361_carry[8]), .S(s2_3_i[7]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_7 ( .A(xo3_r_w_d1r[7]), .B(n1456), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[7]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[8]), .S(dp_cluster_5_s2_3_r[3])
         );
  FA1D0 add_353_U1_6 ( .A(xo4_r_w_d1r[6]), .B(xo6_r_w_d1r[6]), .CI(
        add_353_carry[6]), .CO(add_353_carry[7]), .S(s2_4_r[6]) );
  FA1D0 add_362_U1_6 ( .A(xo4_i_w_d1r[6]), .B(xo6_i_w_d1r[6]), .CI(
        add_362_carry[6]), .CO(add_362_carry[7]), .S(s2_4_i[6]) );
  FA1D0 add_354_U1_7 ( .A(xo5_r_w_d1r[7]), .B(xo7_r_w_d1r[7]), .CI(
        add_354_carry[7]), .CO(add_354_carry[8]), .S(s2_5_r[7]) );
  FA1D0 add_363_U1_7 ( .A(xo5_i_w_d1r[7]), .B(xo7_i_w_d1r[7]), .CI(
        add_363_carry[7]), .CO(add_363_carry[8]), .S(s2_5_i[7]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_5 ( .A(xo7_r_w_d1r[5]), .B(n1590), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[5]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[6]), .S(dp_cluster_4_s2_7_r[5])
         );
  FA1D0 sub_364_U2_5 ( .A(xo4_i_w_d1r[5]), .B(n1664), .CI(sub_364_carry[5]), 
        .CO(sub_364_carry[6]), .S(s2_6_i[5]) );
  FA1D0 sub_365_U2_5 ( .A(xo5_i_w_d1r[5]), .B(n1680), .CI(sub_365_carry[5]), 
        .CO(sub_365_carry[6]), .S(s2_7_i[5]) );
  FA1D0 sub_355_U2_5 ( .A(xo4_r_w_d1r[5]), .B(n1648), .CI(sub_355_carry[5]), 
        .CO(sub_355_carry[6]), .S(s2_6_r[5]) );
  FA1D0 add_349_U1_5 ( .A(xo0_r_w_d1r[5]), .B(xo2_r_w_d1r[5]), .CI(
        add_349_carry[5]), .CO(add_349_carry[6]), .S(s2_0_r[5]) );
  FA1D0 add_358_U1_5 ( .A(xo0_i_w_d1r[5]), .B(xo2_i_w_d1r[5]), .CI(
        add_358_carry[5]), .CO(add_358_carry[6]), .S(s2_0_i[5]) );
  FA1D0 add_350_U1_6 ( .A(xo1_r_w_d1r[6]), .B(xo3_r_w_d1r[6]), .CI(
        add_350_carry[6]), .CO(add_350_carry[7]), .S(s2_1_r[6]) );
  FA1D0 add_359_U1_6 ( .A(xo1_i_w_d1r[6]), .B(xo3_i_w_d1r[6]), .CI(
        add_359_carry[6]), .CO(add_359_carry[7]), .S(s2_1_i[6]) );
  FA1D0 sub_351_U2_5 ( .A(xo0_r_w_d1r[5]), .B(n1520), .CI(sub_351_carry[5]), 
        .CO(sub_351_carry[6]), .S(s2_2_r[5]) );
  FA1D0 sub_360_U2_5 ( .A(xo0_i_w_d1r[5]), .B(n1536), .CI(sub_360_carry[5]), 
        .CO(sub_360_carry[6]), .S(s2_2_i[5]) );
  FA1D0 sub_361_U2_6 ( .A(xo1_i_w_d1r[6]), .B(n1551), .CI(sub_361_carry[6]), 
        .CO(sub_361_carry[7]), .S(s2_3_i[6]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_6 ( .A(xo3_r_w_d1r[6]), .B(n1459), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[6]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[7]), .S(dp_cluster_5_s2_3_r[4])
         );
  FA1D0 add_353_U1_5 ( .A(xo4_r_w_d1r[5]), .B(xo6_r_w_d1r[5]), .CI(
        add_353_carry[5]), .CO(add_353_carry[6]), .S(s2_4_r[5]) );
  FA1D0 add_362_U1_5 ( .A(xo4_i_w_d1r[5]), .B(xo6_i_w_d1r[5]), .CI(
        add_362_carry[5]), .CO(add_362_carry[6]), .S(s2_4_i[5]) );
  FA1D0 add_354_U1_6 ( .A(xo5_r_w_d1r[6]), .B(xo7_r_w_d1r[6]), .CI(
        add_354_carry[6]), .CO(add_354_carry[7]), .S(s2_5_r[6]) );
  FA1D0 add_363_U1_6 ( .A(xo5_i_w_d1r[6]), .B(xo7_i_w_d1r[6]), .CI(
        add_363_carry[6]), .CO(add_363_carry[7]), .S(s2_5_i[6]) );
  FA1D0 sub_334_U2_11 ( .A(xi2_r[58]), .B(n1213), .CI(sub_334_carry[11]), .CO(
        sub_334_carry[12]), .S(s1_6_r[11]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_4 ( .A(xo7_r_w_d1r[4]), .B(n1593), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[4]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[5]), .S(dp_cluster_4_s2_7_r[6])
         );
  FA1D0 sub_364_U2_4 ( .A(xo4_i_w_d1r[4]), .B(n1665), .CI(sub_364_carry[4]), 
        .CO(sub_364_carry[5]), .S(s2_6_i[4]) );
  FA1D0 sub_365_U2_4 ( .A(xo5_i_w_d1r[4]), .B(n1681), .CI(sub_365_carry[4]), 
        .CO(sub_365_carry[5]), .S(s2_7_i[4]) );
  FA1D0 sub_355_U2_4 ( .A(xo4_r_w_d1r[4]), .B(n1649), .CI(sub_355_carry[4]), 
        .CO(sub_355_carry[5]), .S(s2_6_r[4]) );
  FA1D0 add_349_U1_4 ( .A(xo0_r_w_d1r[4]), .B(xo2_r_w_d1r[4]), .CI(
        add_349_carry[4]), .CO(add_349_carry[5]), .S(s2_0_r[4]) );
  FA1D0 add_358_U1_4 ( .A(xo0_i_w_d1r[4]), .B(xo2_i_w_d1r[4]), .CI(
        add_358_carry[4]), .CO(add_358_carry[5]), .S(s2_0_i[4]) );
  FA1D0 add_350_U1_5 ( .A(xo1_r_w_d1r[5]), .B(xo3_r_w_d1r[5]), .CI(
        add_350_carry[5]), .CO(add_350_carry[6]), .S(s2_1_r[5]) );
  FA1D0 add_359_U1_5 ( .A(xo1_i_w_d1r[5]), .B(xo3_i_w_d1r[5]), .CI(
        add_359_carry[5]), .CO(add_359_carry[6]), .S(s2_1_i[5]) );
  FA1D0 sub_351_U2_4 ( .A(xo0_r_w_d1r[4]), .B(n1521), .CI(sub_351_carry[4]), 
        .CO(sub_351_carry[5]), .S(s2_2_r[4]) );
  FA1D0 sub_360_U2_4 ( .A(xo0_i_w_d1r[4]), .B(n1537), .CI(sub_360_carry[4]), 
        .CO(sub_360_carry[5]), .S(s2_2_i[4]) );
  FA1D0 sub_361_U2_5 ( .A(xo1_i_w_d1r[5]), .B(n1552), .CI(sub_361_carry[5]), 
        .CO(sub_361_carry[6]), .S(s2_3_i[5]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_5 ( .A(xo3_r_w_d1r[5]), .B(n1462), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[5]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[6]), .S(dp_cluster_5_s2_3_r[5])
         );
  FA1D0 add_353_U1_4 ( .A(xo4_r_w_d1r[4]), .B(xo6_r_w_d1r[4]), .CI(
        add_353_carry[4]), .CO(add_353_carry[5]), .S(s2_4_r[4]) );
  FA1D0 add_362_U1_4 ( .A(xo4_i_w_d1r[4]), .B(xo6_i_w_d1r[4]), .CI(
        add_362_carry[4]), .CO(add_362_carry[5]), .S(s2_4_i[4]) );
  FA1D0 add_354_U1_5 ( .A(xo5_r_w_d1r[5]), .B(xo7_r_w_d1r[5]), .CI(
        add_354_carry[5]), .CO(add_354_carry[6]), .S(s2_5_r[5]) );
  FA1D0 add_363_U1_5 ( .A(xo5_i_w_d1r[5]), .B(xo7_i_w_d1r[5]), .CI(
        add_363_carry[5]), .CO(add_363_carry[6]), .S(s2_5_i[5]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_3 ( .A(xo7_r_w_d1r[3]), .B(n1596), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[3]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[4]), .S(dp_cluster_4_s2_7_r[7])
         );
  FA1D0 sub_364_U2_3 ( .A(xo4_i_w_d1r[3]), .B(n1666), .CI(sub_364_carry[3]), 
        .CO(sub_364_carry[4]), .S(s2_6_i[3]) );
  FA1D0 sub_355_U2_3 ( .A(xo4_r_w_d1r[3]), .B(n1650), .CI(sub_355_carry[3]), 
        .CO(sub_355_carry[4]), .S(s2_6_r[3]) );
  FA1D0 add_349_U1_3 ( .A(xo0_r_w_d1r[3]), .B(xo2_r_w_d1r[3]), .CI(
        add_349_carry[3]), .CO(add_349_carry[4]), .S(s2_0_r[3]) );
  FA1D0 add_358_U1_3 ( .A(xo0_i_w_d1r[3]), .B(xo2_i_w_d1r[3]), .CI(
        add_358_carry[3]), .CO(add_358_carry[4]), .S(s2_0_i[3]) );
  FA1D0 add_350_U1_4 ( .A(xo1_r_w_d1r[4]), .B(xo3_r_w_d1r[4]), .CI(
        add_350_carry[4]), .CO(add_350_carry[5]), .S(s2_1_r[4]) );
  FA1D0 add_359_U1_4 ( .A(xo1_i_w_d1r[4]), .B(xo3_i_w_d1r[4]), .CI(
        add_359_carry[4]), .CO(add_359_carry[5]), .S(s2_1_i[4]) );
  FA1D0 sub_351_U2_3 ( .A(xo0_r_w_d1r[3]), .B(n1522), .CI(sub_351_carry[3]), 
        .CO(sub_351_carry[4]), .S(s2_2_r[3]) );
  FA1D0 sub_360_U2_3 ( .A(xo0_i_w_d1r[3]), .B(n1538), .CI(sub_360_carry[3]), 
        .CO(sub_360_carry[4]), .S(s2_2_i[3]) );
  FA1D0 sub_361_U2_4 ( .A(xo1_i_w_d1r[4]), .B(n1553), .CI(sub_361_carry[4]), 
        .CO(sub_361_carry[5]), .S(s2_3_i[4]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_4 ( .A(xo3_r_w_d1r[4]), .B(n1465), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[4]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[5]), .S(dp_cluster_5_s2_3_r[6])
         );
  FA1D0 add_353_U1_3 ( .A(xo4_r_w_d1r[3]), .B(xo6_r_w_d1r[3]), .CI(
        add_353_carry[3]), .CO(add_353_carry[4]), .S(s2_4_r[3]) );
  FA1D0 add_362_U1_3 ( .A(xo4_i_w_d1r[3]), .B(xo6_i_w_d1r[3]), .CI(
        add_362_carry[3]), .CO(add_362_carry[4]), .S(s2_4_i[3]) );
  FA1D0 add_354_U1_4 ( .A(xo5_r_w_d1r[4]), .B(xo7_r_w_d1r[4]), .CI(
        add_354_carry[4]), .CO(add_354_carry[5]), .S(s2_5_r[4]) );
  FA1D0 add_363_U1_4 ( .A(xo5_i_w_d1r[4]), .B(xo7_i_w_d1r[4]), .CI(
        add_363_carry[4]), .CO(add_363_carry[5]), .S(s2_5_i[4]) );
  FA1D0 sub_334_U2_10 ( .A(xi2_r[57]), .B(n1214), .CI(sub_334_carry[10]), .CO(
        sub_334_carry[11]), .S(s1_6_r[10]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_2 ( .A(xo7_r_w_d1r[2]), .B(n1599), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[2]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[3]), .S(dp_cluster_4_s2_7_r[8])
         );
  FA1D0 sub_364_U2_2 ( .A(xo4_i_w_d1r[2]), .B(n1667), .CI(sub_364_carry[2]), 
        .CO(sub_364_carry[3]), .S(s2_6_i[2]) );
  FA1D0 sub_365_U2_2 ( .A(xo5_i_w_d1r[2]), .B(n1683), .CI(sub_365_carry[2]), 
        .CO(sub_365_carry[3]), .S(s2_7_i[2]) );
  FA1D0 sub_355_U2_2 ( .A(xo4_r_w_d1r[2]), .B(n1651), .CI(sub_355_carry[2]), 
        .CO(sub_355_carry[3]), .S(s2_6_r[2]) );
  FA1D0 add_349_U1_2 ( .A(xo0_r_w_d1r[2]), .B(xo2_r_w_d1r[2]), .CI(
        add_349_carry[2]), .CO(add_349_carry[3]), .S(s2_0_r[2]) );
  FA1D0 add_358_U1_2 ( .A(xo0_i_w_d1r[2]), .B(xo2_i_w_d1r[2]), .CI(
        add_358_carry[2]), .CO(add_358_carry[3]), .S(s2_0_i[2]) );
  FA1D0 add_350_U1_3 ( .A(xo1_r_w_d1r[3]), .B(xo3_r_w_d1r[3]), .CI(
        add_350_carry[3]), .CO(add_350_carry[4]), .S(s2_1_r[3]) );
  FA1D0 sub_351_U2_2 ( .A(xo0_r_w_d1r[2]), .B(n1523), .CI(sub_351_carry[2]), 
        .CO(sub_351_carry[3]), .S(s2_2_r[2]) );
  FA1D0 sub_360_U2_2 ( .A(xo0_i_w_d1r[2]), .B(n1539), .CI(sub_360_carry[2]), 
        .CO(sub_360_carry[3]), .S(s2_2_i[2]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_3 ( .A(xo3_r_w_d1r[3]), .B(n1468), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[3]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[4]), .S(dp_cluster_5_s2_3_r[7])
         );
  FA1D0 add_353_U1_2 ( .A(xo4_r_w_d1r[2]), .B(xo6_r_w_d1r[2]), .CI(
        add_353_carry[2]), .CO(add_353_carry[3]), .S(s2_4_r[2]) );
  FA1D0 add_362_U1_2 ( .A(xo4_i_w_d1r[2]), .B(xo6_i_w_d1r[2]), .CI(
        add_362_carry[2]), .CO(add_362_carry[3]), .S(s2_4_i[2]) );
  FA1D0 add_354_U1_3 ( .A(xo5_r_w_d1r[3]), .B(xo7_r_w_d1r[3]), .CI(
        add_354_carry[3]), .CO(add_354_carry[4]), .S(s2_5_r[3]) );
  FA1D0 sub_364_U2_1 ( .A(xo4_i_w_d1r[1]), .B(n1668), .CI(sub_364_carry[1]), 
        .CO(sub_364_carry[2]), .S(s2_6_i[1]) );
  FA1D0 sub_355_U2_1 ( .A(xo4_r_w_d1r[1]), .B(n1652), .CI(sub_355_carry[1]), 
        .CO(sub_355_carry[2]), .S(s2_6_r[1]) );
  FA1D0 add_349_U1_1 ( .A(xo0_r_w_d1r[1]), .B(xo2_r_w_d1r[1]), .CI(n918), .CO(
        add_349_carry[2]), .S(s2_0_r[1]) );
  FA1D0 add_358_U1_1 ( .A(xo0_i_w_d1r[1]), .B(xo2_i_w_d1r[1]), .CI(n917), .CO(
        add_358_carry[2]), .S(s2_0_i[1]) );
  FA1D0 add_350_U1_2 ( .A(xo1_r_w_d1r[2]), .B(xo3_r_w_d1r[2]), .CI(
        add_350_carry[2]), .CO(add_350_carry[3]), .S(s2_1_r[2]) );
  FA1D0 add_359_U1_2 ( .A(xo1_i_w_d1r[2]), .B(xo3_i_w_d1r[2]), .CI(
        add_359_carry[2]), .CO(add_359_carry[3]), .S(s2_1_i[2]) );
  FA1D0 sub_351_U2_1 ( .A(xo0_r_w_d1r[1]), .B(n1524), .CI(sub_351_carry[1]), 
        .CO(sub_351_carry[2]), .S(s2_2_r[1]) );
  FA1D0 sub_360_U2_1 ( .A(xo0_i_w_d1r[1]), .B(n1540), .CI(sub_360_carry[1]), 
        .CO(sub_360_carry[2]), .S(s2_2_i[1]) );
  FA1D0 sub_361_U2_2 ( .A(xo1_i_w_d1r[2]), .B(n1555), .CI(sub_361_carry[2]), 
        .CO(sub_361_carry[3]), .S(s2_3_i[2]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_2 ( .A(xo3_r_w_d1r[2]), .B(n1471), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[2]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[3]), .S(dp_cluster_5_s2_3_r[8])
         );
  FA1D0 add_353_U1_1 ( .A(xo4_r_w_d1r[1]), .B(xo6_r_w_d1r[1]), .CI(n916), .CO(
        add_353_carry[2]), .S(s2_4_r[1]) );
  FA1D0 add_362_U1_1 ( .A(xo4_i_w_d1r[1]), .B(xo6_i_w_d1r[1]), .CI(n915), .CO(
        add_362_carry[2]), .S(s2_4_i[1]) );
  FA1D0 add_354_U1_2 ( .A(xo5_r_w_d1r[2]), .B(xo7_r_w_d1r[2]), .CI(
        add_354_carry[2]), .CO(add_354_carry[3]), .S(s2_5_r[2]) );
  FA1D0 add_363_U1_2 ( .A(xo5_i_w_d1r[2]), .B(xo7_i_w_d1r[2]), .CI(
        add_363_carry[2]), .CO(add_363_carry[3]), .S(s2_5_i[2]) );
  FA1D0 sub_334_U2_9 ( .A(xi2_r[56]), .B(n1215), .CI(sub_334_carry[9]), .CO(
        sub_334_carry[10]), .S(s1_6_r[9]) );
  FA1D0 sub_334_U2_8 ( .A(xi2_r[55]), .B(n1216), .CI(sub_334_carry[8]), .CO(
        sub_334_carry[9]), .S(s1_6_r[8]) );
  FA1D0 sub_334_U2_7 ( .A(xi2_r[54]), .B(n1217), .CI(sub_334_carry[7]), .CO(
        sub_334_carry[8]), .S(s1_6_r[7]) );
  FA1D0 sub_334_U2_6 ( .A(xi2_r[53]), .B(n1218), .CI(sub_334_carry[6]), .CO(
        sub_334_carry[7]), .S(s1_6_r[6]) );
  FA1D0 sub_334_U2_5 ( .A(xi2_r[52]), .B(n1219), .CI(sub_334_carry[5]), .CO(
        sub_334_carry[6]), .S(s1_6_r[5]) );
  FA1D0 sub_334_U2_4 ( .A(xi2_r[51]), .B(n1220), .CI(sub_334_carry[4]), .CO(
        sub_334_carry[5]), .S(s1_6_r[4]) );
  FA1D0 sub_334_U2_3 ( .A(xi2_r[50]), .B(n1221), .CI(sub_334_carry[3]), .CO(
        sub_334_carry[4]), .S(s1_6_r[3]) );
  FA1D0 sub_334_U2_2 ( .A(xi2_r[49]), .B(n1222), .CI(sub_334_carry[2]), .CO(
        sub_334_carry[3]), .S(s1_6_r[2]) );
  XOR3D1 sub_365_U2_15 ( .A1(xo5_i_w_d1r[15]), .A2(n1670), .A3(
        sub_365_carry[15]), .Z(s2_7_i[15]) );
  XOR3D1 dp_cluster_4_sub_1_root_sub_444_U2_15 ( .A1(xo7_r_w_d1r[15]), .A2(
        n1560), .A3(dp_cluster_4_sub_1_root_sub_444_carry[15]), .Z(
        dp_cluster_4_s2_7_r[10]) );
  FA1D0 dp_cluster_4_sub_1_root_sub_444_U2_14 ( .A(xo7_r_w_d1r[14]), .B(n1563), 
        .CI(dp_cluster_4_sub_1_root_sub_444_carry[14]), .CO(
        dp_cluster_4_sub_1_root_sub_444_carry[15]), .S(dp_cluster_4_s2_7_r[11]) );
  XOR3D1 add_350_U1_15 ( .A1(xo1_r_w_d1r[15]), .A2(xo3_r_w_d1r[15]), .A3(
        add_350_carry[15]), .Z(s2_1_r[15]) );
  FA1D0 sub_365_U2_14 ( .A(xo5_i_w_d1r[14]), .B(n1671), .CI(sub_365_carry[14]), 
        .CO(sub_365_carry[15]), .S(s2_7_i[14]) );
  XOR3D1 add_359_U1_15 ( .A1(xo1_i_w_d1r[15]), .A2(xo3_i_w_d1r[15]), .A3(
        add_359_carry[15]), .Z(s2_1_i[15]) );
  XOR3D1 sub_361_U2_15 ( .A1(xo1_i_w_d1r[15]), .A2(n1542), .A3(
        sub_361_carry[15]), .Z(s2_3_i[15]) );
  XOR3D1 dp_cluster_5_sub_1_root_sub_440_U2_15 ( .A1(xo3_r_w_d1r[15]), .A2(
        n1432), .A3(dp_cluster_5_sub_1_root_sub_440_carry[15]), .Z(
        dp_cluster_5_s2_3_r[10]) );
  XOR3D1 add_354_U1_15 ( .A1(xo5_r_w_d1r[15]), .A2(xo7_r_w_d1r[15]), .A3(
        add_354_carry[15]), .Z(s2_5_r[15]) );
  FA1D0 add_350_U1_14 ( .A(xo1_r_w_d1r[14]), .B(xo3_r_w_d1r[14]), .CI(
        add_350_carry[14]), .CO(add_350_carry[15]), .S(s2_1_r[14]) );
  XOR3D1 add_363_U1_15 ( .A1(xo5_i_w_d1r[15]), .A2(xo7_i_w_d1r[15]), .A3(
        add_363_carry[15]), .Z(s2_5_i[15]) );
  FA1D0 add_359_U1_14 ( .A(xo1_i_w_d1r[14]), .B(xo3_i_w_d1r[14]), .CI(
        add_359_carry[14]), .CO(add_359_carry[15]), .S(s2_1_i[14]) );
  FA1D0 sub_361_U2_14 ( .A(xo1_i_w_d1r[14]), .B(n1543), .CI(sub_361_carry[14]), 
        .CO(sub_361_carry[15]), .S(s2_3_i[14]) );
  FA1D0 dp_cluster_5_sub_1_root_sub_440_U2_14 ( .A(xo3_r_w_d1r[14]), .B(n1435), 
        .CI(dp_cluster_5_sub_1_root_sub_440_carry[14]), .CO(
        dp_cluster_5_sub_1_root_sub_440_carry[15]), .S(dp_cluster_5_s2_3_r[11]) );
  FA1D0 add_354_U1_14 ( .A(xo5_r_w_d1r[14]), .B(xo7_r_w_d1r[14]), .CI(
        add_354_carry[14]), .CO(add_354_carry[15]), .S(s2_5_r[14]) );
  FA1D0 add_363_U1_14 ( .A(xo5_i_w_d1r[14]), .B(xo7_i_w_d1r[14]), .CI(
        add_363_carry[14]), .CO(add_363_carry[15]), .S(s2_5_i[14]) );
  FA1D0 sub_365_U2_3 ( .A(xo5_i_w_d1r[3]), .B(n1682), .CI(sub_365_carry[3]), 
        .CO(sub_365_carry[4]), .S(s2_7_i[3]) );
  FA1D0 add_359_U1_3 ( .A(xo1_i_w_d1r[3]), .B(xo3_i_w_d1r[3]), .CI(
        add_359_carry[3]), .CO(add_359_carry[4]), .S(s2_1_i[3]) );
  FA1D0 sub_361_U2_3 ( .A(xo1_i_w_d1r[3]), .B(n1554), .CI(sub_361_carry[3]), 
        .CO(sub_361_carry[4]), .S(s2_3_i[3]) );
  FA1D0 add_363_U1_3 ( .A(xo5_i_w_d1r[3]), .B(xo7_i_w_d1r[3]), .CI(
        add_363_carry[3]), .CO(add_363_carry[4]), .S(s2_5_i[3]) );
  XOR3D1 sub_364_U2_15 ( .A1(xo4_i_w_d1r[15]), .A2(n1654), .A3(
        sub_364_carry[15]), .Z(s2_6_i[15]) );
  XOR3D1 sub_355_U2_15 ( .A1(xo4_r_w_d1r[15]), .A2(n1638), .A3(
        sub_355_carry[15]), .Z(s2_6_r[15]) );
  XOR3D1 add_349_U1_15 ( .A1(xo0_r_w_d1r[15]), .A2(xo2_r_w_d1r[15]), .A3(
        add_349_carry[15]), .Z(s2_0_r[15]) );
  XOR3D1 add_358_U1_15 ( .A1(xo0_i_w_d1r[15]), .A2(xo2_i_w_d1r[15]), .A3(
        add_358_carry[15]), .Z(s2_0_i[15]) );
  XOR3D1 sub_351_U2_15 ( .A1(xo0_r_w_d1r[15]), .A2(n1510), .A3(
        sub_351_carry[15]), .Z(s2_2_r[15]) );
  XOR3D1 sub_360_U2_15 ( .A1(xo0_i_w_d1r[15]), .A2(n1526), .A3(
        sub_360_carry[15]), .Z(s2_2_i[15]) );
  XOR3D1 add_353_U1_15 ( .A1(xo4_r_w_d1r[15]), .A2(xo6_r_w_d1r[15]), .A3(
        add_353_carry[15]), .Z(s2_4_r[15]) );
  XOR3D1 add_362_U1_15 ( .A1(xo4_i_w_d1r[15]), .A2(xo6_i_w_d1r[15]), .A3(
        add_362_carry[15]), .Z(s2_4_i[15]) );
  FA1D0 sub_364_U2_14 ( .A(xo4_i_w_d1r[14]), .B(n1655), .CI(sub_364_carry[14]), 
        .CO(sub_364_carry[15]), .S(s2_6_i[14]) );
  FA1D0 sub_355_U2_14 ( .A(xo4_r_w_d1r[14]), .B(n1639), .CI(sub_355_carry[14]), 
        .CO(sub_355_carry[15]), .S(s2_6_r[14]) );
  FA1D0 add_349_U1_14 ( .A(xo0_r_w_d1r[14]), .B(xo2_r_w_d1r[14]), .CI(
        add_349_carry[14]), .CO(add_349_carry[15]), .S(s2_0_r[14]) );
  FA1D0 add_358_U1_14 ( .A(xo0_i_w_d1r[14]), .B(xo2_i_w_d1r[14]), .CI(
        add_358_carry[14]), .CO(add_358_carry[15]), .S(s2_0_i[14]) );
  FA1D0 sub_351_U2_14 ( .A(xo0_r_w_d1r[14]), .B(n1511), .CI(sub_351_carry[14]), 
        .CO(sub_351_carry[15]), .S(s2_2_r[14]) );
  FA1D0 sub_360_U2_14 ( .A(xo0_i_w_d1r[14]), .B(n1527), .CI(sub_360_carry[14]), 
        .CO(sub_360_carry[15]), .S(s2_2_i[14]) );
  FA1D0 add_353_U1_14 ( .A(xo4_r_w_d1r[14]), .B(xo6_r_w_d1r[14]), .CI(
        add_353_carry[14]), .CO(add_353_carry[15]), .S(s2_4_r[14]) );
  FA1D0 add_362_U1_14 ( .A(xo4_i_w_d1r[14]), .B(xo6_i_w_d1r[14]), .CI(
        add_362_carry[14]), .CO(add_362_carry[15]), .S(s2_4_i[14]) );
  FA1D0 sub_342_U2_15 ( .A(xi1_i[62]), .B(n1323), .CI(sub_342_carry[15]), .CO(
        sub_342_carry[16]), .S(s1_5_i[15]) );
  FA1D0 sub_344_U2_15 ( .A(xi3_i[62]), .B(n1355), .CI(sub_344_carry[15]), .CO(
        sub_344_carry[16]), .S(s1_7_i[15]) );
  FA1D0 sub_333_U2_15 ( .A(xi1_r[62]), .B(n1193), .CI(sub_333_carry[15]), .CO(
        sub_333_carry[16]), .S(s1_5_r[15]) );
  FA1D0 sub_342_U2_14 ( .A(xi1_i[61]), .B(n1324), .CI(sub_342_carry[14]), .CO(
        sub_342_carry[15]), .S(s1_5_i[14]) );
  FA1D0 sub_335_U2_15 ( .A(xi3_r[62]), .B(n1225), .CI(sub_335_carry[15]), .CO(
        sub_335_carry[16]), .S(s1_7_r[15]) );
  FA1D0 sub_344_U2_14 ( .A(xi3_i[61]), .B(n1356), .CI(sub_344_carry[14]), .CO(
        sub_344_carry[15]), .S(s1_7_i[14]) );
  FA1D0 sub_333_U2_14 ( .A(xi1_r[61]), .B(n1194), .CI(sub_333_carry[14]), .CO(
        sub_333_carry[15]), .S(s1_5_r[14]) );
  FA1D0 sub_342_U2_13 ( .A(xi1_i[60]), .B(n1325), .CI(sub_342_carry[13]), .CO(
        sub_342_carry[14]), .S(s1_5_i[13]) );
  FA1D0 sub_335_U2_14 ( .A(xi3_r[61]), .B(n1226), .CI(sub_335_carry[14]), .CO(
        sub_335_carry[15]), .S(s1_7_r[14]) );
  FA1D0 sub_344_U2_13 ( .A(xi3_i[60]), .B(n1357), .CI(sub_344_carry[13]), .CO(
        sub_344_carry[14]), .S(s1_7_i[13]) );
  FA1D0 sub_333_U2_13 ( .A(xi1_r[60]), .B(n1195), .CI(sub_333_carry[13]), .CO(
        sub_333_carry[14]), .S(s1_5_r[13]) );
  FA1D0 sub_342_U2_12 ( .A(xi1_i[59]), .B(n1326), .CI(sub_342_carry[12]), .CO(
        sub_342_carry[13]), .S(s1_5_i[12]) );
  FA1D0 sub_335_U2_13 ( .A(xi3_r[60]), .B(n1227), .CI(sub_335_carry[13]), .CO(
        sub_335_carry[14]), .S(s1_7_r[13]) );
  FA1D0 sub_344_U2_12 ( .A(xi3_i[59]), .B(n1358), .CI(sub_344_carry[12]), .CO(
        sub_344_carry[13]), .S(s1_7_i[12]) );
  FA1D0 sub_333_U2_12 ( .A(xi1_r[59]), .B(n1196), .CI(sub_333_carry[12]), .CO(
        sub_333_carry[13]), .S(s1_5_r[12]) );
  FA1D0 sub_342_U2_11 ( .A(xi1_i[58]), .B(n1327), .CI(sub_342_carry[11]), .CO(
        sub_342_carry[12]), .S(s1_5_i[11]) );
  FA1D0 sub_335_U2_12 ( .A(xi3_r[59]), .B(n1228), .CI(sub_335_carry[12]), .CO(
        sub_335_carry[13]), .S(s1_7_r[12]) );
  FA1D0 sub_344_U2_11 ( .A(xi3_i[58]), .B(n1359), .CI(sub_344_carry[11]), .CO(
        sub_344_carry[12]), .S(s1_7_i[11]) );
  FA1D0 sub_333_U2_11 ( .A(xi1_r[58]), .B(n1197), .CI(sub_333_carry[11]), .CO(
        sub_333_carry[12]), .S(s1_5_r[11]) );
  FA1D0 sub_342_U2_10 ( .A(xi1_i[57]), .B(n1328), .CI(sub_342_carry[10]), .CO(
        sub_342_carry[11]), .S(s1_5_i[10]) );
  FA1D0 sub_335_U2_11 ( .A(xi3_r[58]), .B(n1229), .CI(sub_335_carry[11]), .CO(
        sub_335_carry[12]), .S(s1_7_r[11]) );
  FA1D0 sub_344_U2_10 ( .A(xi3_i[57]), .B(n1360), .CI(sub_344_carry[10]), .CO(
        sub_344_carry[11]), .S(s1_7_i[10]) );
  FA1D0 sub_333_U2_10 ( .A(xi1_r[57]), .B(n1198), .CI(sub_333_carry[10]), .CO(
        sub_333_carry[11]), .S(s1_5_r[10]) );
  FA1D0 sub_342_U2_9 ( .A(xi1_i[56]), .B(n1329), .CI(sub_342_carry[9]), .CO(
        sub_342_carry[10]), .S(s1_5_i[9]) );
  FA1D0 sub_335_U2_10 ( .A(xi3_r[57]), .B(n1230), .CI(sub_335_carry[10]), .CO(
        sub_335_carry[11]), .S(s1_7_r[10]) );
  FA1D0 sub_344_U2_9 ( .A(xi3_i[56]), .B(n1361), .CI(sub_344_carry[9]), .CO(
        sub_344_carry[10]), .S(s1_7_i[9]) );
  FA1D0 sub_333_U2_9 ( .A(xi1_r[56]), .B(n1199), .CI(sub_333_carry[9]), .CO(
        sub_333_carry[10]), .S(s1_5_r[9]) );
  FA1D0 sub_342_U2_8 ( .A(xi1_i[55]), .B(n1330), .CI(sub_342_carry[8]), .CO(
        sub_342_carry[9]), .S(s1_5_i[8]) );
  FA1D0 sub_335_U2_9 ( .A(xi3_r[56]), .B(n1231), .CI(sub_335_carry[9]), .CO(
        sub_335_carry[10]), .S(s1_7_r[9]) );
  FA1D0 sub_344_U2_8 ( .A(xi3_i[55]), .B(n1362), .CI(sub_344_carry[8]), .CO(
        sub_344_carry[9]), .S(s1_7_i[8]) );
  FA1D0 sub_333_U2_8 ( .A(xi1_r[55]), .B(n1200), .CI(sub_333_carry[8]), .CO(
        sub_333_carry[9]), .S(s1_5_r[8]) );
  FA1D0 sub_342_U2_7 ( .A(xi1_i[54]), .B(n1331), .CI(sub_342_carry[7]), .CO(
        sub_342_carry[8]), .S(s1_5_i[7]) );
  FA1D0 sub_335_U2_8 ( .A(xi3_r[55]), .B(n1232), .CI(sub_335_carry[8]), .CO(
        sub_335_carry[9]), .S(s1_7_r[8]) );
  FA1D0 sub_344_U2_7 ( .A(xi3_i[54]), .B(n1363), .CI(sub_344_carry[7]), .CO(
        sub_344_carry[8]), .S(s1_7_i[7]) );
  FA1D0 sub_333_U2_7 ( .A(xi1_r[54]), .B(n1201), .CI(sub_333_carry[7]), .CO(
        sub_333_carry[8]), .S(s1_5_r[7]) );
  FA1D0 sub_335_U2_7 ( .A(xi3_r[54]), .B(n1233), .CI(sub_335_carry[7]), .CO(
        sub_335_carry[8]), .S(s1_7_r[7]) );
  FA1D0 sub_333_U2_6 ( .A(xi1_r[53]), .B(n1202), .CI(sub_333_carry[6]), .CO(
        sub_333_carry[7]), .S(s1_5_r[6]) );
  FA1D0 sub_342_U2_6 ( .A(xi1_i[53]), .B(n1332), .CI(sub_342_carry[6]), .CO(
        sub_342_carry[7]), .S(s1_5_i[6]) );
  FA1D0 sub_335_U2_6 ( .A(xi3_r[53]), .B(n1234), .CI(sub_335_carry[6]), .CO(
        sub_335_carry[7]), .S(s1_7_r[6]) );
  FA1D0 sub_344_U2_6 ( .A(xi3_i[53]), .B(n1364), .CI(sub_344_carry[6]), .CO(
        sub_344_carry[7]), .S(s1_7_i[6]) );
  FA1D0 sub_333_U2_5 ( .A(xi1_r[52]), .B(n1203), .CI(sub_333_carry[5]), .CO(
        sub_333_carry[6]), .S(s1_5_r[5]) );
  FA1D0 sub_333_U2_1 ( .A(xi1_r[48]), .B(n1207), .CI(sub_333_carry[1]), .CO(
        sub_333_carry[2]), .S(s1_5_r[1]) );
  FA1D0 sub_342_U2_5 ( .A(xi1_i[52]), .B(n1333), .CI(sub_342_carry[5]), .CO(
        sub_342_carry[6]), .S(s1_5_i[5]) );
  FA1D0 sub_342_U2_1 ( .A(xi1_i[48]), .B(n1337), .CI(sub_342_carry[1]), .CO(
        sub_342_carry[2]), .S(s1_5_i[1]) );
  FA1D0 sub_335_U2_5 ( .A(xi3_r[52]), .B(n1235), .CI(sub_335_carry[5]), .CO(
        sub_335_carry[6]), .S(s1_7_r[5]) );
  FA1D0 sub_335_U2_1 ( .A(xi3_r[48]), .B(n1239), .CI(sub_335_carry[1]), .CO(
        sub_335_carry[2]), .S(s1_7_r[1]) );
  FA1D0 sub_344_U2_5 ( .A(xi3_i[52]), .B(n1365), .CI(sub_344_carry[5]), .CO(
        sub_344_carry[6]), .S(s1_7_i[5]) );
  FA1D0 sub_344_U2_1 ( .A(xi3_i[48]), .B(n1369), .CI(sub_344_carry[1]), .CO(
        sub_344_carry[2]), .S(s1_7_i[1]) );
  FA1D0 sub_333_U2_4 ( .A(xi1_r[51]), .B(n1204), .CI(sub_333_carry[4]), .CO(
        sub_333_carry[5]), .S(s1_5_r[4]) );
  FA1D0 sub_342_U2_4 ( .A(xi1_i[51]), .B(n1334), .CI(sub_342_carry[4]), .CO(
        sub_342_carry[5]), .S(s1_5_i[4]) );
  FA1D0 sub_335_U2_4 ( .A(xi3_r[51]), .B(n1236), .CI(sub_335_carry[4]), .CO(
        sub_335_carry[5]), .S(s1_7_r[4]) );
  FA1D0 sub_344_U2_4 ( .A(xi3_i[51]), .B(n1366), .CI(sub_344_carry[4]), .CO(
        sub_344_carry[5]), .S(s1_7_i[4]) );
  FA1D0 sub_333_U2_3 ( .A(xi1_r[50]), .B(n1205), .CI(sub_333_carry[3]), .CO(
        sub_333_carry[4]), .S(s1_5_r[3]) );
  FA1D0 sub_342_U2_3 ( .A(xi1_i[50]), .B(n1335), .CI(sub_342_carry[3]), .CO(
        sub_342_carry[4]), .S(s1_5_i[3]) );
  FA1D0 sub_335_U2_3 ( .A(xi3_r[50]), .B(n1237), .CI(sub_335_carry[3]), .CO(
        sub_335_carry[4]), .S(s1_7_r[3]) );
  FA1D0 sub_344_U2_3 ( .A(xi3_i[50]), .B(n1367), .CI(sub_344_carry[3]), .CO(
        sub_344_carry[4]), .S(s1_7_i[3]) );
  FA1D0 sub_342_U2_2 ( .A(xi1_i[49]), .B(n1336), .CI(sub_342_carry[2]), .CO(
        sub_342_carry[3]), .S(s1_5_i[2]) );
  FA1D0 sub_344_U2_2 ( .A(xi3_i[49]), .B(n1368), .CI(sub_344_carry[2]), .CO(
        sub_344_carry[3]), .S(s1_7_i[2]) );
  FA1D0 sub_333_U2_2 ( .A(xi1_r[49]), .B(n1206), .CI(sub_333_carry[2]), .CO(
        sub_333_carry[3]), .S(s1_5_r[2]) );
  FA1D0 sub_335_U2_2 ( .A(xi3_r[49]), .B(n1238), .CI(sub_335_carry[2]), .CO(
        sub_335_carry[3]), .S(s1_7_r[2]) );
  XOR3D1 sub_333_U2_16 ( .A1(xi1_r[63]), .A2(n1192), .A3(sub_333_carry[16]), 
        .Z(s1_5_r[16]) );
  XOR3D1 sub_335_U2_16 ( .A1(xi3_r[63]), .A2(n1224), .A3(sub_335_carry[16]), 
        .Z(s1_7_r[16]) );
  XOR3D1 sub_342_U2_16 ( .A1(xi1_i[63]), .A2(n1322), .A3(sub_342_carry[16]), 
        .Z(s1_5_i[16]) );
  XOR3D1 sub_344_U2_16 ( .A1(xi3_i[63]), .A2(n1354), .A3(sub_344_carry[16]), 
        .Z(s1_7_i[16]) );
  FA1D0 sub_385_U2_2 ( .A(s2_6_i[2]), .B(n1598), .CI(sub_385_carry[2]), .CO(
        sub_385_carry[3]), .S(s3_7_i[2]) );
  FA1D0 sub_385_U2_3 ( .A(s2_6_i[3]), .B(n1595), .CI(sub_385_carry[3]), .CO(
        sub_385_carry[4]), .S(s3_7_i[3]) );
  FA1D0 sub_385_U2_4 ( .A(s2_6_i[4]), .B(n1592), .CI(sub_385_carry[4]), .CO(
        sub_385_carry[5]), .S(s3_7_i[4]) );
  FA1D0 sub_385_U2_5 ( .A(s2_6_i[5]), .B(n1589), .CI(sub_385_carry[5]), .CO(
        sub_385_carry[6]), .S(s3_7_i[5]) );
  FA1D0 sub_385_U2_6 ( .A(s2_6_i[6]), .B(n1586), .CI(sub_385_carry[6]), .CO(
        sub_385_carry[7]), .S(s3_7_i[6]) );
  FA1D0 sub_385_U2_7 ( .A(s2_6_i[7]), .B(n1583), .CI(sub_385_carry[7]), .CO(
        sub_385_carry[8]), .S(s3_7_i[7]) );
  FA1D0 sub_381_U2_7 ( .A(s2_2_i[7]), .B(n1455), .CI(sub_381_carry[7]), .CO(
        sub_381_carry[8]), .S(s3_3_i[7]) );
  FA1D0 sub_381_U2_6 ( .A(s2_2_i[6]), .B(n1458), .CI(sub_381_carry[6]), .CO(
        sub_381_carry[7]), .S(s3_3_i[6]) );
  FA1D0 sub_381_U2_5 ( .A(s2_2_i[5]), .B(n1461), .CI(sub_381_carry[5]), .CO(
        sub_381_carry[6]), .S(s3_3_i[5]) );
  FA1D0 sub_381_U2_4 ( .A(s2_2_i[4]), .B(n1464), .CI(sub_381_carry[4]), .CO(
        sub_381_carry[5]), .S(s3_3_i[4]) );
  FA1D0 sub_381_U2_3 ( .A(s2_2_i[3]), .B(n1467), .CI(sub_381_carry[3]), .CO(
        sub_381_carry[4]), .S(s3_3_i[3]) );
  FA1D0 sub_381_U2_2 ( .A(s2_2_i[2]), .B(n1470), .CI(sub_381_carry[2]), .CO(
        sub_381_carry[3]), .S(s3_3_i[2]) );
  XOR3D1 sub_385_U2_15 ( .A1(s2_6_i[15]), .A2(n1559), .A3(sub_385_carry[15]), 
        .Z(s3_7_i[15]) );
  XOR3D1 sub_376_U2_15 ( .A1(s2_6_r[15]), .A2(n1607), .A3(sub_376_carry[15]), 
        .Z(s3_7_r[15]) );
  XOR3D1 add_369_U1_15 ( .A1(s2_0_r[15]), .A2(s2_1_r[15]), .A3(
        add_369_carry[15]), .Z(s3_0_r[15]) );
  XOR3D1 add_378_U1_15 ( .A1(s2_0_i[15]), .A2(s2_1_i[15]), .A3(
        add_378_carry[15]), .Z(s3_0_i[15]) );
  XOR3D1 sub_370_U2_15 ( .A1(s2_0_r[15]), .A2(n1430), .A3(sub_370_carry[15]), 
        .Z(s3_1_r[15]) );
  XOR3D1 sub_379_U2_15 ( .A1(s2_0_i[15]), .A2(n1478), .A3(sub_379_carry[15]), 
        .Z(s3_1_i[15]) );
  XOR3D1 add_371_U1_15 ( .A1(s2_2_r[15]), .A2(s2_3_i[15]), .A3(
        add_371_carry[15]), .Z(s3_2_r[15]) );
  XOR3D1 add_380_U1_15 ( .A1(s2_2_i[15]), .A2(dp_cluster_5_s2_3_r[10]), .A3(
        add_380_carry[15]), .Z(s3_2_i[15]) );
  XOR3D1 sub_372_U2_15 ( .A1(s2_2_r[15]), .A2(n1479), .A3(sub_372_carry[15]), 
        .Z(s3_3_r[15]) );
  XOR3D1 sub_381_U2_15 ( .A1(s2_2_i[15]), .A2(n1431), .A3(sub_381_carry[15]), 
        .Z(s3_3_i[15]) );
  XOR3D1 add_373_U1_15 ( .A1(s2_4_r[15]), .A2(s2_5_r[15]), .A3(
        add_373_carry[15]), .Z(s3_4_r[15]) );
  XOR3D1 add_382_U1_15 ( .A1(s2_4_i[15]), .A2(s2_5_i[15]), .A3(
        add_382_carry[15]), .Z(s3_4_i[15]) );
  XOR3D1 sub_374_U2_15 ( .A1(s2_4_r[15]), .A2(n1558), .A3(sub_374_carry[15]), 
        .Z(s3_5_r[15]) );
  XOR3D1 sub_383_U2_15 ( .A1(s2_4_i[15]), .A2(n1606), .A3(sub_383_carry[15]), 
        .Z(s3_5_i[15]) );
  XOR3D1 add_375_U1_15 ( .A1(s2_6_r[15]), .A2(s2_7_i[15]), .A3(
        add_375_carry[15]), .Z(s3_6_r[15]) );
  XOR3D1 add_384_U1_15 ( .A1(s2_6_i[15]), .A2(dp_cluster_4_s2_7_r[10]), .A3(
        add_384_carry[15]), .Z(s3_6_i[15]) );
  FA1D0 sub_385_U2_1 ( .A(s2_6_i[1]), .B(n1601), .CI(sub_385_carry[1]), .CO(
        sub_385_carry[2]), .S(s3_7_i[1]) );
  FA1D0 sub_385_U2_8 ( .A(s2_6_i[8]), .B(n1580), .CI(sub_385_carry[8]), .CO(
        sub_385_carry[9]), .S(s3_7_i[8]) );
  FA1D0 sub_385_U2_9 ( .A(s2_6_i[9]), .B(n1577), .CI(sub_385_carry[9]), .CO(
        sub_385_carry[10]), .S(s3_7_i[9]) );
  FA1D0 sub_385_U2_10 ( .A(s2_6_i[10]), .B(n1574), .CI(sub_385_carry[10]), 
        .CO(sub_385_carry[11]), .S(s3_7_i[10]) );
  FA1D0 sub_385_U2_11 ( .A(s2_6_i[11]), .B(n1571), .CI(sub_385_carry[11]), 
        .CO(sub_385_carry[12]), .S(s3_7_i[11]) );
  FA1D0 sub_385_U2_12 ( .A(s2_6_i[12]), .B(n1568), .CI(sub_385_carry[12]), 
        .CO(sub_385_carry[13]), .S(s3_7_i[12]) );
  FA1D0 sub_385_U2_13 ( .A(s2_6_i[13]), .B(n1565), .CI(sub_385_carry[13]), 
        .CO(sub_385_carry[14]), .S(s3_7_i[13]) );
  FA1D0 sub_385_U2_14 ( .A(s2_6_i[14]), .B(n1562), .CI(sub_385_carry[14]), 
        .CO(sub_385_carry[15]), .S(s3_7_i[14]) );
  FA1D0 sub_376_U2_1 ( .A(s2_6_r[1]), .B(n1635), .CI(sub_376_carry[1]), .CO(
        sub_376_carry[2]), .S(s3_7_r[1]) );
  FA1D0 sub_376_U2_2 ( .A(s2_6_r[2]), .B(n1633), .CI(sub_376_carry[2]), .CO(
        sub_376_carry[3]), .S(s3_7_r[2]) );
  FA1D0 sub_376_U2_3 ( .A(s2_6_r[3]), .B(n1631), .CI(sub_376_carry[3]), .CO(
        sub_376_carry[4]), .S(s3_7_r[3]) );
  FA1D0 sub_376_U2_4 ( .A(s2_6_r[4]), .B(n1629), .CI(sub_376_carry[4]), .CO(
        sub_376_carry[5]), .S(s3_7_r[4]) );
  FA1D0 sub_376_U2_5 ( .A(s2_6_r[5]), .B(n1627), .CI(sub_376_carry[5]), .CO(
        sub_376_carry[6]), .S(s3_7_r[5]) );
  FA1D0 sub_376_U2_6 ( .A(s2_6_r[6]), .B(n1625), .CI(sub_376_carry[6]), .CO(
        sub_376_carry[7]), .S(s3_7_r[6]) );
  FA1D0 sub_376_U2_7 ( .A(s2_6_r[7]), .B(n1623), .CI(sub_376_carry[7]), .CO(
        sub_376_carry[8]), .S(s3_7_r[7]) );
  FA1D0 sub_376_U2_8 ( .A(s2_6_r[8]), .B(n1621), .CI(sub_376_carry[8]), .CO(
        sub_376_carry[9]), .S(s3_7_r[8]) );
  FA1D0 sub_376_U2_9 ( .A(s2_6_r[9]), .B(n1619), .CI(sub_376_carry[9]), .CO(
        sub_376_carry[10]), .S(s3_7_r[9]) );
  FA1D0 sub_376_U2_10 ( .A(s2_6_r[10]), .B(n1617), .CI(sub_376_carry[10]), 
        .CO(sub_376_carry[11]), .S(s3_7_r[10]) );
  FA1D0 sub_376_U2_11 ( .A(s2_6_r[11]), .B(n1615), .CI(sub_376_carry[11]), 
        .CO(sub_376_carry[12]), .S(s3_7_r[11]) );
  FA1D0 sub_376_U2_12 ( .A(s2_6_r[12]), .B(n1613), .CI(sub_376_carry[12]), 
        .CO(sub_376_carry[13]), .S(s3_7_r[12]) );
  FA1D0 sub_376_U2_13 ( .A(s2_6_r[13]), .B(n1611), .CI(sub_376_carry[13]), 
        .CO(sub_376_carry[14]), .S(s3_7_r[13]) );
  FA1D0 sub_376_U2_14 ( .A(s2_6_r[14]), .B(n1609), .CI(sub_376_carry[14]), 
        .CO(sub_376_carry[15]), .S(s3_7_r[14]) );
  FA1D0 add_369_U1_14 ( .A(s2_0_r[14]), .B(s2_1_r[14]), .CI(add_369_carry[14]), 
        .CO(add_369_carry[15]), .S(s3_0_r[14]) );
  FA1D0 add_369_U1_13 ( .A(s2_0_r[13]), .B(s2_1_r[13]), .CI(add_369_carry[13]), 
        .CO(add_369_carry[14]), .S(s3_0_r[13]) );
  FA1D0 add_369_U1_12 ( .A(s2_0_r[12]), .B(s2_1_r[12]), .CI(add_369_carry[12]), 
        .CO(add_369_carry[13]), .S(s3_0_r[12]) );
  FA1D0 add_369_U1_11 ( .A(s2_0_r[11]), .B(s2_1_r[11]), .CI(add_369_carry[11]), 
        .CO(add_369_carry[12]), .S(s3_0_r[11]) );
  FA1D0 add_369_U1_10 ( .A(s2_0_r[10]), .B(s2_1_r[10]), .CI(add_369_carry[10]), 
        .CO(add_369_carry[11]), .S(s3_0_r[10]) );
  FA1D0 add_369_U1_9 ( .A(s2_0_r[9]), .B(s2_1_r[9]), .CI(add_369_carry[9]), 
        .CO(add_369_carry[10]), .S(s3_0_r[9]) );
  FA1D0 add_369_U1_8 ( .A(s2_0_r[8]), .B(s2_1_r[8]), .CI(add_369_carry[8]), 
        .CO(add_369_carry[9]), .S(s3_0_r[8]) );
  FA1D0 add_369_U1_7 ( .A(s2_0_r[7]), .B(s2_1_r[7]), .CI(add_369_carry[7]), 
        .CO(add_369_carry[8]), .S(s3_0_r[7]) );
  FA1D0 add_369_U1_6 ( .A(s2_0_r[6]), .B(s2_1_r[6]), .CI(add_369_carry[6]), 
        .CO(add_369_carry[7]), .S(s3_0_r[6]) );
  FA1D0 add_369_U1_5 ( .A(s2_0_r[5]), .B(s2_1_r[5]), .CI(add_369_carry[5]), 
        .CO(add_369_carry[6]), .S(s3_0_r[5]) );
  FA1D0 add_369_U1_4 ( .A(s2_0_r[4]), .B(s2_1_r[4]), .CI(add_369_carry[4]), 
        .CO(add_369_carry[5]), .S(s3_0_r[4]) );
  FA1D0 add_369_U1_3 ( .A(s2_0_r[3]), .B(s2_1_r[3]), .CI(add_369_carry[3]), 
        .CO(add_369_carry[4]), .S(s3_0_r[3]) );
  FA1D0 add_369_U1_2 ( .A(s2_0_r[2]), .B(s2_1_r[2]), .CI(add_369_carry[2]), 
        .CO(add_369_carry[3]), .S(s3_0_r[2]) );
  FA1D0 add_369_U1_1 ( .A(s2_0_r[1]), .B(s2_1_r[1]), .CI(n910), .CO(
        add_369_carry[2]), .S(s3_0_r[1]) );
  FA1D0 add_378_U1_14 ( .A(s2_0_i[14]), .B(s2_1_i[14]), .CI(add_378_carry[14]), 
        .CO(add_378_carry[15]), .S(s3_0_i[14]) );
  FA1D0 add_378_U1_13 ( .A(s2_0_i[13]), .B(s2_1_i[13]), .CI(add_378_carry[13]), 
        .CO(add_378_carry[14]), .S(s3_0_i[13]) );
  FA1D0 add_378_U1_12 ( .A(s2_0_i[12]), .B(s2_1_i[12]), .CI(add_378_carry[12]), 
        .CO(add_378_carry[13]), .S(s3_0_i[12]) );
  FA1D0 add_378_U1_11 ( .A(s2_0_i[11]), .B(s2_1_i[11]), .CI(add_378_carry[11]), 
        .CO(add_378_carry[12]), .S(s3_0_i[11]) );
  FA1D0 add_378_U1_10 ( .A(s2_0_i[10]), .B(s2_1_i[10]), .CI(add_378_carry[10]), 
        .CO(add_378_carry[11]), .S(s3_0_i[10]) );
  FA1D0 add_378_U1_9 ( .A(s2_0_i[9]), .B(s2_1_i[9]), .CI(add_378_carry[9]), 
        .CO(add_378_carry[10]), .S(s3_0_i[9]) );
  FA1D0 add_378_U1_8 ( .A(s2_0_i[8]), .B(s2_1_i[8]), .CI(add_378_carry[8]), 
        .CO(add_378_carry[9]), .S(s3_0_i[8]) );
  FA1D0 add_378_U1_7 ( .A(s2_0_i[7]), .B(s2_1_i[7]), .CI(add_378_carry[7]), 
        .CO(add_378_carry[8]), .S(s3_0_i[7]) );
  FA1D0 add_378_U1_6 ( .A(s2_0_i[6]), .B(s2_1_i[6]), .CI(add_378_carry[6]), 
        .CO(add_378_carry[7]), .S(s3_0_i[6]) );
  FA1D0 add_378_U1_5 ( .A(s2_0_i[5]), .B(s2_1_i[5]), .CI(add_378_carry[5]), 
        .CO(add_378_carry[6]), .S(s3_0_i[5]) );
  FA1D0 add_378_U1_4 ( .A(s2_0_i[4]), .B(s2_1_i[4]), .CI(add_378_carry[4]), 
        .CO(add_378_carry[5]), .S(s3_0_i[4]) );
  FA1D0 add_378_U1_3 ( .A(s2_0_i[3]), .B(s2_1_i[3]), .CI(add_378_carry[3]), 
        .CO(add_378_carry[4]), .S(s3_0_i[3]) );
  FA1D0 add_378_U1_2 ( .A(s2_0_i[2]), .B(s2_1_i[2]), .CI(add_378_carry[2]), 
        .CO(add_378_carry[3]), .S(s3_0_i[2]) );
  FA1D0 add_378_U1_1 ( .A(s2_0_i[1]), .B(s2_1_i[1]), .CI(n909), .CO(
        add_378_carry[2]), .S(s3_0_i[1]) );
  FA1D0 sub_370_U2_14 ( .A(s2_0_r[14]), .B(n1433), .CI(sub_370_carry[14]), 
        .CO(sub_370_carry[15]), .S(s3_1_r[14]) );
  FA1D0 sub_370_U2_13 ( .A(s2_0_r[13]), .B(n1436), .CI(sub_370_carry[13]), 
        .CO(sub_370_carry[14]), .S(s3_1_r[13]) );
  FA1D0 sub_370_U2_12 ( .A(s2_0_r[12]), .B(n1439), .CI(sub_370_carry[12]), 
        .CO(sub_370_carry[13]), .S(s3_1_r[12]) );
  FA1D0 sub_370_U2_11 ( .A(s2_0_r[11]), .B(n1442), .CI(sub_370_carry[11]), 
        .CO(sub_370_carry[12]), .S(s3_1_r[11]) );
  FA1D0 sub_370_U2_10 ( .A(s2_0_r[10]), .B(n1445), .CI(sub_370_carry[10]), 
        .CO(sub_370_carry[11]), .S(s3_1_r[10]) );
  FA1D0 sub_370_U2_9 ( .A(s2_0_r[9]), .B(n1448), .CI(sub_370_carry[9]), .CO(
        sub_370_carry[10]), .S(s3_1_r[9]) );
  FA1D0 sub_370_U2_8 ( .A(s2_0_r[8]), .B(n1451), .CI(sub_370_carry[8]), .CO(
        sub_370_carry[9]), .S(s3_1_r[8]) );
  FA1D0 sub_370_U2_7 ( .A(s2_0_r[7]), .B(n1454), .CI(sub_370_carry[7]), .CO(
        sub_370_carry[8]), .S(s3_1_r[7]) );
  FA1D0 sub_370_U2_6 ( .A(s2_0_r[6]), .B(n1457), .CI(sub_370_carry[6]), .CO(
        sub_370_carry[7]), .S(s3_1_r[6]) );
  FA1D0 sub_370_U2_5 ( .A(s2_0_r[5]), .B(n1460), .CI(sub_370_carry[5]), .CO(
        sub_370_carry[6]), .S(s3_1_r[5]) );
  FA1D0 sub_370_U2_4 ( .A(s2_0_r[4]), .B(n1463), .CI(sub_370_carry[4]), .CO(
        sub_370_carry[5]), .S(s3_1_r[4]) );
  FA1D0 sub_370_U2_3 ( .A(s2_0_r[3]), .B(n1466), .CI(sub_370_carry[3]), .CO(
        sub_370_carry[4]), .S(s3_1_r[3]) );
  FA1D0 sub_370_U2_2 ( .A(s2_0_r[2]), .B(n1469), .CI(sub_370_carry[2]), .CO(
        sub_370_carry[3]), .S(s3_1_r[2]) );
  FA1D0 sub_370_U2_1 ( .A(s2_0_r[1]), .B(n1472), .CI(sub_370_carry[1]), .CO(
        sub_370_carry[2]), .S(s3_1_r[1]) );
  FA1D0 sub_379_U2_14 ( .A(s2_0_i[14]), .B(n1480), .CI(sub_379_carry[14]), 
        .CO(sub_379_carry[15]), .S(s3_1_i[14]) );
  FA1D0 sub_379_U2_13 ( .A(s2_0_i[13]), .B(n1482), .CI(sub_379_carry[13]), 
        .CO(sub_379_carry[14]), .S(s3_1_i[13]) );
  FA1D0 sub_379_U2_12 ( .A(s2_0_i[12]), .B(n1484), .CI(sub_379_carry[12]), 
        .CO(sub_379_carry[13]), .S(s3_1_i[12]) );
  FA1D0 sub_379_U2_11 ( .A(s2_0_i[11]), .B(n1486), .CI(sub_379_carry[11]), 
        .CO(sub_379_carry[12]), .S(s3_1_i[11]) );
  FA1D0 sub_379_U2_10 ( .A(s2_0_i[10]), .B(n1488), .CI(sub_379_carry[10]), 
        .CO(sub_379_carry[11]), .S(s3_1_i[10]) );
  FA1D0 sub_379_U2_9 ( .A(s2_0_i[9]), .B(n1490), .CI(sub_379_carry[9]), .CO(
        sub_379_carry[10]), .S(s3_1_i[9]) );
  FA1D0 sub_379_U2_8 ( .A(s2_0_i[8]), .B(n1492), .CI(sub_379_carry[8]), .CO(
        sub_379_carry[9]), .S(s3_1_i[8]) );
  FA1D0 sub_379_U2_7 ( .A(s2_0_i[7]), .B(n1494), .CI(sub_379_carry[7]), .CO(
        sub_379_carry[8]), .S(s3_1_i[7]) );
  FA1D0 sub_379_U2_6 ( .A(s2_0_i[6]), .B(n1496), .CI(sub_379_carry[6]), .CO(
        sub_379_carry[7]), .S(s3_1_i[6]) );
  FA1D0 sub_379_U2_5 ( .A(s2_0_i[5]), .B(n1498), .CI(sub_379_carry[5]), .CO(
        sub_379_carry[6]), .S(s3_1_i[5]) );
  FA1D0 sub_379_U2_4 ( .A(s2_0_i[4]), .B(n1500), .CI(sub_379_carry[4]), .CO(
        sub_379_carry[5]), .S(s3_1_i[4]) );
  FA1D0 sub_379_U2_3 ( .A(s2_0_i[3]), .B(n1502), .CI(sub_379_carry[3]), .CO(
        sub_379_carry[4]), .S(s3_1_i[3]) );
  FA1D0 sub_379_U2_2 ( .A(s2_0_i[2]), .B(n1504), .CI(sub_379_carry[2]), .CO(
        sub_379_carry[3]), .S(s3_1_i[2]) );
  FA1D0 sub_379_U2_1 ( .A(s2_0_i[1]), .B(n1506), .CI(sub_379_carry[1]), .CO(
        sub_379_carry[2]), .S(s3_1_i[1]) );
  FA1D0 add_371_U1_14 ( .A(s2_2_r[14]), .B(s2_3_i[14]), .CI(add_371_carry[14]), 
        .CO(add_371_carry[15]), .S(s3_2_r[14]) );
  FA1D0 add_371_U1_13 ( .A(s2_2_r[13]), .B(s2_3_i[13]), .CI(add_371_carry[13]), 
        .CO(add_371_carry[14]), .S(s3_2_r[13]) );
  FA1D0 add_371_U1_12 ( .A(s2_2_r[12]), .B(s2_3_i[12]), .CI(add_371_carry[12]), 
        .CO(add_371_carry[13]), .S(s3_2_r[12]) );
  FA1D0 add_371_U1_11 ( .A(s2_2_r[11]), .B(s2_3_i[11]), .CI(add_371_carry[11]), 
        .CO(add_371_carry[12]), .S(s3_2_r[11]) );
  FA1D0 add_371_U1_10 ( .A(s2_2_r[10]), .B(s2_3_i[10]), .CI(add_371_carry[10]), 
        .CO(add_371_carry[11]), .S(s3_2_r[10]) );
  FA1D0 add_371_U1_9 ( .A(s2_2_r[9]), .B(s2_3_i[9]), .CI(add_371_carry[9]), 
        .CO(add_371_carry[10]), .S(s3_2_r[9]) );
  FA1D0 add_371_U1_8 ( .A(s2_2_r[8]), .B(s2_3_i[8]), .CI(add_371_carry[8]), 
        .CO(add_371_carry[9]), .S(s3_2_r[8]) );
  FA1D0 add_371_U1_7 ( .A(s2_2_r[7]), .B(s2_3_i[7]), .CI(add_371_carry[7]), 
        .CO(add_371_carry[8]), .S(s3_2_r[7]) );
  FA1D0 add_371_U1_6 ( .A(s2_2_r[6]), .B(s2_3_i[6]), .CI(add_371_carry[6]), 
        .CO(add_371_carry[7]), .S(s3_2_r[6]) );
  FA1D0 add_371_U1_5 ( .A(s2_2_r[5]), .B(s2_3_i[5]), .CI(add_371_carry[5]), 
        .CO(add_371_carry[6]), .S(s3_2_r[5]) );
  FA1D0 add_371_U1_4 ( .A(s2_2_r[4]), .B(s2_3_i[4]), .CI(add_371_carry[4]), 
        .CO(add_371_carry[5]), .S(s3_2_r[4]) );
  FA1D0 add_371_U1_3 ( .A(s2_2_r[3]), .B(s2_3_i[3]), .CI(add_371_carry[3]), 
        .CO(add_371_carry[4]), .S(s3_2_r[3]) );
  FA1D0 add_371_U1_2 ( .A(s2_2_r[2]), .B(s2_3_i[2]), .CI(add_371_carry[2]), 
        .CO(add_371_carry[3]), .S(s3_2_r[2]) );
  FA1D0 add_371_U1_1 ( .A(s2_2_r[1]), .B(s2_3_i[1]), .CI(n914), .CO(
        add_371_carry[2]), .S(s3_2_r[1]) );
  FA1D0 add_380_U1_14 ( .A(s2_2_i[14]), .B(dp_cluster_5_s2_3_r[11]), .CI(
        add_380_carry[14]), .CO(add_380_carry[15]), .S(s3_2_i[14]) );
  FA1D0 add_380_U1_13 ( .A(s2_2_i[13]), .B(dp_cluster_5_s2_3_r[12]), .CI(
        add_380_carry[13]), .CO(add_380_carry[14]), .S(s3_2_i[13]) );
  FA1D0 add_380_U1_12 ( .A(s2_2_i[12]), .B(dp_cluster_5_s2_3_r[13]), .CI(
        add_380_carry[12]), .CO(add_380_carry[13]), .S(s3_2_i[12]) );
  FA1D0 add_380_U1_11 ( .A(s2_2_i[11]), .B(dp_cluster_5_s2_3_r[14]), .CI(
        add_380_carry[11]), .CO(add_380_carry[12]), .S(s3_2_i[11]) );
  FA1D0 add_380_U1_10 ( .A(s2_2_i[10]), .B(dp_cluster_5_s2_3_r[15]), .CI(
        add_380_carry[10]), .CO(add_380_carry[11]), .S(s3_2_i[10]) );
  FA1D0 add_380_U1_9 ( .A(s2_2_i[9]), .B(dp_cluster_5_s2_3_r[1]), .CI(
        add_380_carry[9]), .CO(add_380_carry[10]), .S(s3_2_i[9]) );
  FA1D0 add_380_U1_8 ( .A(s2_2_i[8]), .B(dp_cluster_5_s2_3_r[2]), .CI(
        add_380_carry[8]), .CO(add_380_carry[9]), .S(s3_2_i[8]) );
  FA1D0 add_380_U1_7 ( .A(s2_2_i[7]), .B(dp_cluster_5_s2_3_r[3]), .CI(
        add_380_carry[7]), .CO(add_380_carry[8]), .S(s3_2_i[7]) );
  FA1D0 add_380_U1_6 ( .A(s2_2_i[6]), .B(dp_cluster_5_s2_3_r[4]), .CI(
        add_380_carry[6]), .CO(add_380_carry[7]), .S(s3_2_i[6]) );
  FA1D0 add_380_U1_5 ( .A(s2_2_i[5]), .B(dp_cluster_5_s2_3_r[5]), .CI(
        add_380_carry[5]), .CO(add_380_carry[6]), .S(s3_2_i[5]) );
  FA1D0 add_380_U1_4 ( .A(s2_2_i[4]), .B(dp_cluster_5_s2_3_r[6]), .CI(
        add_380_carry[4]), .CO(add_380_carry[5]), .S(s3_2_i[4]) );
  FA1D0 add_380_U1_3 ( .A(s2_2_i[3]), .B(dp_cluster_5_s2_3_r[7]), .CI(
        add_380_carry[3]), .CO(add_380_carry[4]), .S(s3_2_i[3]) );
  FA1D0 add_380_U1_2 ( .A(s2_2_i[2]), .B(dp_cluster_5_s2_3_r[8]), .CI(
        add_380_carry[2]), .CO(add_380_carry[3]), .S(s3_2_i[2]) );
  FA1D0 add_380_U1_1 ( .A(s2_2_i[1]), .B(dp_cluster_5_s2_3_r[9]), .CI(n913), 
        .CO(add_380_carry[2]), .S(s3_2_i[1]) );
  FA1D0 sub_372_U2_14 ( .A(s2_2_r[14]), .B(n1481), .CI(sub_372_carry[14]), 
        .CO(sub_372_carry[15]), .S(s3_3_r[14]) );
  FA1D0 sub_372_U2_13 ( .A(s2_2_r[13]), .B(n1483), .CI(sub_372_carry[13]), 
        .CO(sub_372_carry[14]), .S(s3_3_r[13]) );
  FA1D0 sub_372_U2_12 ( .A(s2_2_r[12]), .B(n1485), .CI(sub_372_carry[12]), 
        .CO(sub_372_carry[13]), .S(s3_3_r[12]) );
  FA1D0 sub_372_U2_11 ( .A(s2_2_r[11]), .B(n1487), .CI(sub_372_carry[11]), 
        .CO(sub_372_carry[12]), .S(s3_3_r[11]) );
  FA1D0 sub_372_U2_10 ( .A(s2_2_r[10]), .B(n1489), .CI(sub_372_carry[10]), 
        .CO(sub_372_carry[11]), .S(s3_3_r[10]) );
  FA1D0 sub_372_U2_9 ( .A(s2_2_r[9]), .B(n1491), .CI(sub_372_carry[9]), .CO(
        sub_372_carry[10]), .S(s3_3_r[9]) );
  FA1D0 sub_372_U2_8 ( .A(s2_2_r[8]), .B(n1493), .CI(sub_372_carry[8]), .CO(
        sub_372_carry[9]), .S(s3_3_r[8]) );
  FA1D0 sub_372_U2_7 ( .A(s2_2_r[7]), .B(n1495), .CI(sub_372_carry[7]), .CO(
        sub_372_carry[8]), .S(s3_3_r[7]) );
  FA1D0 sub_372_U2_6 ( .A(s2_2_r[6]), .B(n1497), .CI(sub_372_carry[6]), .CO(
        sub_372_carry[7]), .S(s3_3_r[6]) );
  FA1D0 sub_372_U2_5 ( .A(s2_2_r[5]), .B(n1499), .CI(sub_372_carry[5]), .CO(
        sub_372_carry[6]), .S(s3_3_r[5]) );
  FA1D0 sub_372_U2_4 ( .A(s2_2_r[4]), .B(n1501), .CI(sub_372_carry[4]), .CO(
        sub_372_carry[5]), .S(s3_3_r[4]) );
  FA1D0 sub_372_U2_3 ( .A(s2_2_r[3]), .B(n1503), .CI(sub_372_carry[3]), .CO(
        sub_372_carry[4]), .S(s3_3_r[3]) );
  FA1D0 sub_372_U2_2 ( .A(s2_2_r[2]), .B(n1505), .CI(sub_372_carry[2]), .CO(
        sub_372_carry[3]), .S(s3_3_r[2]) );
  FA1D0 sub_372_U2_1 ( .A(s2_2_r[1]), .B(n1507), .CI(sub_372_carry[1]), .CO(
        sub_372_carry[2]), .S(s3_3_r[1]) );
  FA1D0 sub_381_U2_14 ( .A(s2_2_i[14]), .B(n1434), .CI(sub_381_carry[14]), 
        .CO(sub_381_carry[15]), .S(s3_3_i[14]) );
  FA1D0 sub_381_U2_13 ( .A(s2_2_i[13]), .B(n1437), .CI(sub_381_carry[13]), 
        .CO(sub_381_carry[14]), .S(s3_3_i[13]) );
  FA1D0 sub_381_U2_12 ( .A(s2_2_i[12]), .B(n1440), .CI(sub_381_carry[12]), 
        .CO(sub_381_carry[13]), .S(s3_3_i[12]) );
  FA1D0 sub_381_U2_11 ( .A(s2_2_i[11]), .B(n1443), .CI(sub_381_carry[11]), 
        .CO(sub_381_carry[12]), .S(s3_3_i[11]) );
  FA1D0 sub_381_U2_10 ( .A(s2_2_i[10]), .B(n1446), .CI(sub_381_carry[10]), 
        .CO(sub_381_carry[11]), .S(s3_3_i[10]) );
  FA1D0 sub_381_U2_9 ( .A(s2_2_i[9]), .B(n1449), .CI(sub_381_carry[9]), .CO(
        sub_381_carry[10]), .S(s3_3_i[9]) );
  FA1D0 sub_381_U2_8 ( .A(s2_2_i[8]), .B(n1452), .CI(sub_381_carry[8]), .CO(
        sub_381_carry[9]), .S(s3_3_i[8]) );
  FA1D0 sub_381_U2_1 ( .A(s2_2_i[1]), .B(n1473), .CI(sub_381_carry[1]), .CO(
        sub_381_carry[2]), .S(s3_3_i[1]) );
  FA1D0 add_373_U1_14 ( .A(s2_4_r[14]), .B(s2_5_r[14]), .CI(add_373_carry[14]), 
        .CO(add_373_carry[15]), .S(s3_4_r[14]) );
  FA1D0 add_373_U1_13 ( .A(s2_4_r[13]), .B(s2_5_r[13]), .CI(add_373_carry[13]), 
        .CO(add_373_carry[14]), .S(s3_4_r[13]) );
  FA1D0 add_373_U1_12 ( .A(s2_4_r[12]), .B(s2_5_r[12]), .CI(add_373_carry[12]), 
        .CO(add_373_carry[13]), .S(s3_4_r[12]) );
  FA1D0 add_373_U1_11 ( .A(s2_4_r[11]), .B(s2_5_r[11]), .CI(add_373_carry[11]), 
        .CO(add_373_carry[12]), .S(s3_4_r[11]) );
  FA1D0 add_373_U1_10 ( .A(s2_4_r[10]), .B(s2_5_r[10]), .CI(add_373_carry[10]), 
        .CO(add_373_carry[11]), .S(s3_4_r[10]) );
  FA1D0 add_373_U1_9 ( .A(s2_4_r[9]), .B(s2_5_r[9]), .CI(add_373_carry[9]), 
        .CO(add_373_carry[10]), .S(s3_4_r[9]) );
  FA1D0 add_373_U1_8 ( .A(s2_4_r[8]), .B(s2_5_r[8]), .CI(add_373_carry[8]), 
        .CO(add_373_carry[9]), .S(s3_4_r[8]) );
  FA1D0 add_373_U1_7 ( .A(s2_4_r[7]), .B(s2_5_r[7]), .CI(add_373_carry[7]), 
        .CO(add_373_carry[8]), .S(s3_4_r[7]) );
  FA1D0 add_373_U1_6 ( .A(s2_4_r[6]), .B(s2_5_r[6]), .CI(add_373_carry[6]), 
        .CO(add_373_carry[7]), .S(s3_4_r[6]) );
  FA1D0 add_373_U1_5 ( .A(s2_4_r[5]), .B(s2_5_r[5]), .CI(add_373_carry[5]), 
        .CO(add_373_carry[6]), .S(s3_4_r[5]) );
  FA1D0 add_373_U1_4 ( .A(s2_4_r[4]), .B(s2_5_r[4]), .CI(add_373_carry[4]), 
        .CO(add_373_carry[5]), .S(s3_4_r[4]) );
  FA1D0 add_373_U1_3 ( .A(s2_4_r[3]), .B(s2_5_r[3]), .CI(add_373_carry[3]), 
        .CO(add_373_carry[4]), .S(s3_4_r[3]) );
  FA1D0 add_373_U1_2 ( .A(s2_4_r[2]), .B(s2_5_r[2]), .CI(add_373_carry[2]), 
        .CO(add_373_carry[3]), .S(s3_4_r[2]) );
  FA1D0 add_373_U1_1 ( .A(s2_4_r[1]), .B(s2_5_r[1]), .CI(n908), .CO(
        add_373_carry[2]), .S(s3_4_r[1]) );
  FA1D0 add_382_U1_14 ( .A(s2_4_i[14]), .B(s2_5_i[14]), .CI(add_382_carry[14]), 
        .CO(add_382_carry[15]), .S(s3_4_i[14]) );
  FA1D0 add_382_U1_13 ( .A(s2_4_i[13]), .B(s2_5_i[13]), .CI(add_382_carry[13]), 
        .CO(add_382_carry[14]), .S(s3_4_i[13]) );
  FA1D0 add_382_U1_12 ( .A(s2_4_i[12]), .B(s2_5_i[12]), .CI(add_382_carry[12]), 
        .CO(add_382_carry[13]), .S(s3_4_i[12]) );
  FA1D0 add_382_U1_11 ( .A(s2_4_i[11]), .B(s2_5_i[11]), .CI(add_382_carry[11]), 
        .CO(add_382_carry[12]), .S(s3_4_i[11]) );
  FA1D0 add_382_U1_10 ( .A(s2_4_i[10]), .B(s2_5_i[10]), .CI(add_382_carry[10]), 
        .CO(add_382_carry[11]), .S(s3_4_i[10]) );
  FA1D0 add_382_U1_9 ( .A(s2_4_i[9]), .B(s2_5_i[9]), .CI(add_382_carry[9]), 
        .CO(add_382_carry[10]), .S(s3_4_i[9]) );
  FA1D0 add_382_U1_8 ( .A(s2_4_i[8]), .B(s2_5_i[8]), .CI(add_382_carry[8]), 
        .CO(add_382_carry[9]), .S(s3_4_i[8]) );
  FA1D0 add_382_U1_7 ( .A(s2_4_i[7]), .B(s2_5_i[7]), .CI(add_382_carry[7]), 
        .CO(add_382_carry[8]), .S(s3_4_i[7]) );
  FA1D0 add_382_U1_6 ( .A(s2_4_i[6]), .B(s2_5_i[6]), .CI(add_382_carry[6]), 
        .CO(add_382_carry[7]), .S(s3_4_i[6]) );
  FA1D0 add_382_U1_5 ( .A(s2_4_i[5]), .B(s2_5_i[5]), .CI(add_382_carry[5]), 
        .CO(add_382_carry[6]), .S(s3_4_i[5]) );
  FA1D0 add_382_U1_4 ( .A(s2_4_i[4]), .B(s2_5_i[4]), .CI(add_382_carry[4]), 
        .CO(add_382_carry[5]), .S(s3_4_i[4]) );
  FA1D0 add_382_U1_3 ( .A(s2_4_i[3]), .B(s2_5_i[3]), .CI(add_382_carry[3]), 
        .CO(add_382_carry[4]), .S(s3_4_i[3]) );
  FA1D0 add_382_U1_2 ( .A(s2_4_i[2]), .B(s2_5_i[2]), .CI(add_382_carry[2]), 
        .CO(add_382_carry[3]), .S(s3_4_i[2]) );
  FA1D0 add_382_U1_1 ( .A(s2_4_i[1]), .B(s2_5_i[1]), .CI(n907), .CO(
        add_382_carry[2]), .S(s3_4_i[1]) );
  FA1D0 sub_374_U2_14 ( .A(s2_4_r[14]), .B(n1561), .CI(sub_374_carry[14]), 
        .CO(sub_374_carry[15]), .S(s3_5_r[14]) );
  FA1D0 sub_374_U2_13 ( .A(s2_4_r[13]), .B(n1564), .CI(sub_374_carry[13]), 
        .CO(sub_374_carry[14]), .S(s3_5_r[13]) );
  FA1D0 sub_374_U2_12 ( .A(s2_4_r[12]), .B(n1567), .CI(sub_374_carry[12]), 
        .CO(sub_374_carry[13]), .S(s3_5_r[12]) );
  FA1D0 sub_374_U2_11 ( .A(s2_4_r[11]), .B(n1570), .CI(sub_374_carry[11]), 
        .CO(sub_374_carry[12]), .S(s3_5_r[11]) );
  FA1D0 sub_374_U2_10 ( .A(s2_4_r[10]), .B(n1573), .CI(sub_374_carry[10]), 
        .CO(sub_374_carry[11]), .S(s3_5_r[10]) );
  FA1D0 sub_374_U2_9 ( .A(s2_4_r[9]), .B(n1576), .CI(sub_374_carry[9]), .CO(
        sub_374_carry[10]), .S(s3_5_r[9]) );
  FA1D0 sub_374_U2_8 ( .A(s2_4_r[8]), .B(n1579), .CI(sub_374_carry[8]), .CO(
        sub_374_carry[9]), .S(s3_5_r[8]) );
  FA1D0 sub_374_U2_7 ( .A(s2_4_r[7]), .B(n1582), .CI(sub_374_carry[7]), .CO(
        sub_374_carry[8]), .S(s3_5_r[7]) );
  FA1D0 sub_374_U2_6 ( .A(s2_4_r[6]), .B(n1585), .CI(sub_374_carry[6]), .CO(
        sub_374_carry[7]), .S(s3_5_r[6]) );
  FA1D0 sub_374_U2_5 ( .A(s2_4_r[5]), .B(n1588), .CI(sub_374_carry[5]), .CO(
        sub_374_carry[6]), .S(s3_5_r[5]) );
  FA1D0 sub_374_U2_4 ( .A(s2_4_r[4]), .B(n1591), .CI(sub_374_carry[4]), .CO(
        sub_374_carry[5]), .S(s3_5_r[4]) );
  FA1D0 sub_374_U2_3 ( .A(s2_4_r[3]), .B(n1594), .CI(sub_374_carry[3]), .CO(
        sub_374_carry[4]), .S(s3_5_r[3]) );
  FA1D0 sub_374_U2_2 ( .A(s2_4_r[2]), .B(n1597), .CI(sub_374_carry[2]), .CO(
        sub_374_carry[3]), .S(s3_5_r[2]) );
  FA1D0 sub_374_U2_1 ( .A(s2_4_r[1]), .B(n1600), .CI(sub_374_carry[1]), .CO(
        sub_374_carry[2]), .S(s3_5_r[1]) );
  FA1D0 sub_383_U2_14 ( .A(s2_4_i[14]), .B(n1608), .CI(sub_383_carry[14]), 
        .CO(sub_383_carry[15]), .S(s3_5_i[14]) );
  FA1D0 sub_383_U2_13 ( .A(s2_4_i[13]), .B(n1610), .CI(sub_383_carry[13]), 
        .CO(sub_383_carry[14]), .S(s3_5_i[13]) );
  FA1D0 sub_383_U2_12 ( .A(s2_4_i[12]), .B(n1612), .CI(sub_383_carry[12]), 
        .CO(sub_383_carry[13]), .S(s3_5_i[12]) );
  FA1D0 sub_383_U2_11 ( .A(s2_4_i[11]), .B(n1614), .CI(sub_383_carry[11]), 
        .CO(sub_383_carry[12]), .S(s3_5_i[11]) );
  FA1D0 sub_383_U2_10 ( .A(s2_4_i[10]), .B(n1616), .CI(sub_383_carry[10]), 
        .CO(sub_383_carry[11]), .S(s3_5_i[10]) );
  FA1D0 sub_383_U2_9 ( .A(s2_4_i[9]), .B(n1618), .CI(sub_383_carry[9]), .CO(
        sub_383_carry[10]), .S(s3_5_i[9]) );
  FA1D0 sub_383_U2_8 ( .A(s2_4_i[8]), .B(n1620), .CI(sub_383_carry[8]), .CO(
        sub_383_carry[9]), .S(s3_5_i[8]) );
  FA1D0 sub_383_U2_7 ( .A(s2_4_i[7]), .B(n1622), .CI(sub_383_carry[7]), .CO(
        sub_383_carry[8]), .S(s3_5_i[7]) );
  FA1D0 sub_383_U2_6 ( .A(s2_4_i[6]), .B(n1624), .CI(sub_383_carry[6]), .CO(
        sub_383_carry[7]), .S(s3_5_i[6]) );
  FA1D0 sub_383_U2_5 ( .A(s2_4_i[5]), .B(n1626), .CI(sub_383_carry[5]), .CO(
        sub_383_carry[6]), .S(s3_5_i[5]) );
  FA1D0 sub_383_U2_4 ( .A(s2_4_i[4]), .B(n1628), .CI(sub_383_carry[4]), .CO(
        sub_383_carry[5]), .S(s3_5_i[4]) );
  FA1D0 sub_383_U2_3 ( .A(s2_4_i[3]), .B(n1630), .CI(sub_383_carry[3]), .CO(
        sub_383_carry[4]), .S(s3_5_i[3]) );
  FA1D0 sub_383_U2_2 ( .A(s2_4_i[2]), .B(n1632), .CI(sub_383_carry[2]), .CO(
        sub_383_carry[3]), .S(s3_5_i[2]) );
  FA1D0 sub_383_U2_1 ( .A(s2_4_i[1]), .B(n1634), .CI(sub_383_carry[1]), .CO(
        sub_383_carry[2]), .S(s3_5_i[1]) );
  FA1D0 add_375_U1_14 ( .A(s2_6_r[14]), .B(s2_7_i[14]), .CI(add_375_carry[14]), 
        .CO(add_375_carry[15]), .S(s3_6_r[14]) );
  FA1D0 add_375_U1_13 ( .A(s2_6_r[13]), .B(s2_7_i[13]), .CI(add_375_carry[13]), 
        .CO(add_375_carry[14]), .S(s3_6_r[13]) );
  FA1D0 add_375_U1_12 ( .A(s2_6_r[12]), .B(s2_7_i[12]), .CI(add_375_carry[12]), 
        .CO(add_375_carry[13]), .S(s3_6_r[12]) );
  FA1D0 add_375_U1_11 ( .A(s2_6_r[11]), .B(s2_7_i[11]), .CI(add_375_carry[11]), 
        .CO(add_375_carry[12]), .S(s3_6_r[11]) );
  FA1D0 add_375_U1_10 ( .A(s2_6_r[10]), .B(s2_7_i[10]), .CI(add_375_carry[10]), 
        .CO(add_375_carry[11]), .S(s3_6_r[10]) );
  FA1D0 add_375_U1_9 ( .A(s2_6_r[9]), .B(s2_7_i[9]), .CI(add_375_carry[9]), 
        .CO(add_375_carry[10]), .S(s3_6_r[9]) );
  FA1D0 add_375_U1_8 ( .A(s2_6_r[8]), .B(s2_7_i[8]), .CI(add_375_carry[8]), 
        .CO(add_375_carry[9]), .S(s3_6_r[8]) );
  FA1D0 add_375_U1_7 ( .A(s2_6_r[7]), .B(s2_7_i[7]), .CI(add_375_carry[7]), 
        .CO(add_375_carry[8]), .S(s3_6_r[7]) );
  FA1D0 add_375_U1_6 ( .A(s2_6_r[6]), .B(s2_7_i[6]), .CI(add_375_carry[6]), 
        .CO(add_375_carry[7]), .S(s3_6_r[6]) );
  FA1D0 add_375_U1_5 ( .A(s2_6_r[5]), .B(s2_7_i[5]), .CI(add_375_carry[5]), 
        .CO(add_375_carry[6]), .S(s3_6_r[5]) );
  FA1D0 add_375_U1_4 ( .A(s2_6_r[4]), .B(s2_7_i[4]), .CI(add_375_carry[4]), 
        .CO(add_375_carry[5]), .S(s3_6_r[4]) );
  FA1D0 add_375_U1_3 ( .A(s2_6_r[3]), .B(s2_7_i[3]), .CI(add_375_carry[3]), 
        .CO(add_375_carry[4]), .S(s3_6_r[3]) );
  FA1D0 add_375_U1_2 ( .A(s2_6_r[2]), .B(s2_7_i[2]), .CI(add_375_carry[2]), 
        .CO(add_375_carry[3]), .S(s3_6_r[2]) );
  FA1D0 add_375_U1_1 ( .A(s2_6_r[1]), .B(s2_7_i[1]), .CI(n912), .CO(
        add_375_carry[2]), .S(s3_6_r[1]) );
  FA1D0 add_384_U1_14 ( .A(s2_6_i[14]), .B(dp_cluster_4_s2_7_r[11]), .CI(
        add_384_carry[14]), .CO(add_384_carry[15]), .S(s3_6_i[14]) );
  FA1D0 add_384_U1_13 ( .A(s2_6_i[13]), .B(dp_cluster_4_s2_7_r[12]), .CI(
        add_384_carry[13]), .CO(add_384_carry[14]), .S(s3_6_i[13]) );
  FA1D0 add_384_U1_12 ( .A(s2_6_i[12]), .B(dp_cluster_4_s2_7_r[13]), .CI(
        add_384_carry[12]), .CO(add_384_carry[13]), .S(s3_6_i[12]) );
  FA1D0 add_384_U1_11 ( .A(s2_6_i[11]), .B(dp_cluster_4_s2_7_r[14]), .CI(
        add_384_carry[11]), .CO(add_384_carry[12]), .S(s3_6_i[11]) );
  FA1D0 add_384_U1_10 ( .A(s2_6_i[10]), .B(dp_cluster_4_s2_7_r[15]), .CI(
        add_384_carry[10]), .CO(add_384_carry[11]), .S(s3_6_i[10]) );
  FA1D0 add_384_U1_9 ( .A(s2_6_i[9]), .B(dp_cluster_4_s2_7_r[1]), .CI(
        add_384_carry[9]), .CO(add_384_carry[10]), .S(s3_6_i[9]) );
  FA1D0 add_384_U1_8 ( .A(s2_6_i[8]), .B(dp_cluster_4_s2_7_r[2]), .CI(
        add_384_carry[8]), .CO(add_384_carry[9]), .S(s3_6_i[8]) );
  FA1D0 add_384_U1_7 ( .A(s2_6_i[7]), .B(dp_cluster_4_s2_7_r[3]), .CI(
        add_384_carry[7]), .CO(add_384_carry[8]), .S(s3_6_i[7]) );
  FA1D0 add_384_U1_6 ( .A(s2_6_i[6]), .B(dp_cluster_4_s2_7_r[4]), .CI(
        add_384_carry[6]), .CO(add_384_carry[7]), .S(s3_6_i[6]) );
  FA1D0 add_384_U1_5 ( .A(s2_6_i[5]), .B(dp_cluster_4_s2_7_r[5]), .CI(
        add_384_carry[5]), .CO(add_384_carry[6]), .S(s3_6_i[5]) );
  FA1D0 add_384_U1_4 ( .A(s2_6_i[4]), .B(dp_cluster_4_s2_7_r[6]), .CI(
        add_384_carry[4]), .CO(add_384_carry[5]), .S(s3_6_i[4]) );
  FA1D0 add_384_U1_3 ( .A(s2_6_i[3]), .B(dp_cluster_4_s2_7_r[7]), .CI(
        add_384_carry[3]), .CO(add_384_carry[4]), .S(s3_6_i[3]) );
  FA1D0 add_384_U1_2 ( .A(s2_6_i[2]), .B(dp_cluster_4_s2_7_r[8]), .CI(
        add_384_carry[2]), .CO(add_384_carry[3]), .S(s3_6_i[2]) );
  FA1D0 add_384_U1_1 ( .A(s2_6_i[1]), .B(dp_cluster_4_s2_7_r[9]), .CI(n911), 
        .CO(add_384_carry[2]), .S(s3_6_i[1]) );
  XOR3D1 dp_cluster_2_sub_487_C409_U2_27 ( .A1(dp_cluster_2_N28), .A2(n906), 
        .A3(dp_cluster_2_sub_487_C409_carry[27]), .Z(s1_5_tmp_r[15]) );
  XOR3D1 dp_cluster_0_sub_487_C412_U2_27 ( .A1(dp_cluster_0_N84), .A2(n905), 
        .A3(dp_cluster_0_sub_487_C412_carry[27]), .Z(s1_7_tmp_r[15]) );
  XOR3D1 dp_cluster_3_add_514_C415_U1_27 ( .A1(dp_cluster_3_N140), .A2(
        dp_cluster_3_N168), .A3(dp_cluster_3_add_514_C415_carry[27]), .Z(
        s1_5_tmp_i[15]) );
  XOR3D1 dp_cluster_1_add_514_C418_U1_27 ( .A1(dp_cluster_1_N196), .A2(
        dp_cluster_1_N224), .A3(dp_cluster_1_add_514_C418_carry[27]), .Z(
        s1_7_tmp_i[15]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_26 ( .A(dp_cluster_2_N27), .B(n1240), 
        .CI(dp_cluster_2_sub_487_C409_carry[26]), .CO(
        dp_cluster_2_sub_487_C409_carry[27]), .S(s1_5_tmp_r[14]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_26 ( .A(dp_cluster_0_N83), .B(n1273), 
        .CI(dp_cluster_0_sub_487_C412_carry[26]), .CO(
        dp_cluster_0_sub_487_C412_carry[27]), .S(s1_7_tmp_r[14]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_12 ( .A(dp_cluster_2_N13), .B(n1256), 
        .CI(dp_cluster_2_sub_487_C409_carry[12]), .CO(
        dp_cluster_2_sub_487_C409_carry[13]), .S(s1_5_tmp_r[0]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_26 ( .A(dp_cluster_3_N139), .B(
        dp_cluster_3_N167), .CI(dp_cluster_3_add_514_C415_carry[26]), .CO(
        dp_cluster_3_add_514_C415_carry[27]), .S(s1_5_tmp_i[14]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_12 ( .A(dp_cluster_3_N125), .B(
        dp_cluster_3_N153), .CI(dp_cluster_3_add_514_C415_carry[12]), .CO(
        dp_cluster_3_add_514_C415_carry[13]), .S(s1_5_tmp_i[0]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_12 ( .A(dp_cluster_0_N69), .B(n1289), 
        .CI(dp_cluster_0_sub_487_C412_carry[12]), .CO(
        dp_cluster_0_sub_487_C412_carry[13]), .S(s1_7_tmp_r[0]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_26 ( .A(dp_cluster_1_N195), .B(
        dp_cluster_1_N223), .CI(dp_cluster_1_add_514_C418_carry[26]), .CO(
        dp_cluster_1_add_514_C418_carry[27]), .S(s1_7_tmp_i[14]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_12 ( .A(dp_cluster_1_N181), .B(
        dp_cluster_1_N209), .CI(dp_cluster_1_add_514_C418_carry[12]), .CO(
        dp_cluster_1_add_514_C418_carry[13]), .S(s1_7_tmp_i[0]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_25 ( .A(dp_cluster_2_N26), .B(n1241), 
        .CI(dp_cluster_2_sub_487_C409_carry[25]), .CO(
        dp_cluster_2_sub_487_C409_carry[26]), .S(s1_5_tmp_r[13]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_24 ( .A(dp_cluster_2_N25), .B(n1242), 
        .CI(dp_cluster_2_sub_487_C409_carry[24]), .CO(
        dp_cluster_2_sub_487_C409_carry[25]), .S(s1_5_tmp_r[12]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_23 ( .A(dp_cluster_2_N24), .B(n1243), 
        .CI(dp_cluster_2_sub_487_C409_carry[23]), .CO(
        dp_cluster_2_sub_487_C409_carry[24]), .S(s1_5_tmp_r[11]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_22 ( .A(dp_cluster_2_N23), .B(n1244), 
        .CI(dp_cluster_2_sub_487_C409_carry[22]), .CO(
        dp_cluster_2_sub_487_C409_carry[23]), .S(s1_5_tmp_r[10]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_21 ( .A(dp_cluster_2_N22), .B(n1245), 
        .CI(dp_cluster_2_sub_487_C409_carry[21]), .CO(
        dp_cluster_2_sub_487_C409_carry[22]), .S(s1_5_tmp_r[9]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_20 ( .A(dp_cluster_2_N21), .B(n1246), 
        .CI(dp_cluster_2_sub_487_C409_carry[20]), .CO(
        dp_cluster_2_sub_487_C409_carry[21]), .S(s1_5_tmp_r[8]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_19 ( .A(dp_cluster_2_N20), .B(n1247), 
        .CI(dp_cluster_2_sub_487_C409_carry[19]), .CO(
        dp_cluster_2_sub_487_C409_carry[20]), .S(s1_5_tmp_r[7]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_18 ( .A(dp_cluster_2_N19), .B(n1248), 
        .CI(dp_cluster_2_sub_487_C409_carry[18]), .CO(
        dp_cluster_2_sub_487_C409_carry[19]), .S(s1_5_tmp_r[6]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_17 ( .A(dp_cluster_2_N18), .B(n1249), 
        .CI(dp_cluster_2_sub_487_C409_carry[17]), .CO(
        dp_cluster_2_sub_487_C409_carry[18]), .S(s1_5_tmp_r[5]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_16 ( .A(dp_cluster_2_N17), .B(n1250), 
        .CI(dp_cluster_2_sub_487_C409_carry[16]), .CO(
        dp_cluster_2_sub_487_C409_carry[17]), .S(s1_5_tmp_r[4]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_25 ( .A(dp_cluster_0_N82), .B(n1274), 
        .CI(dp_cluster_0_sub_487_C412_carry[25]), .CO(
        dp_cluster_0_sub_487_C412_carry[26]), .S(s1_7_tmp_r[13]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_24 ( .A(dp_cluster_0_N81), .B(n1275), 
        .CI(dp_cluster_0_sub_487_C412_carry[24]), .CO(
        dp_cluster_0_sub_487_C412_carry[25]), .S(s1_7_tmp_r[12]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_23 ( .A(dp_cluster_0_N80), .B(n1276), 
        .CI(dp_cluster_0_sub_487_C412_carry[23]), .CO(
        dp_cluster_0_sub_487_C412_carry[24]), .S(s1_7_tmp_r[11]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_22 ( .A(dp_cluster_0_N79), .B(n1277), 
        .CI(dp_cluster_0_sub_487_C412_carry[22]), .CO(
        dp_cluster_0_sub_487_C412_carry[23]), .S(s1_7_tmp_r[10]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_21 ( .A(dp_cluster_0_N78), .B(n1278), 
        .CI(dp_cluster_0_sub_487_C412_carry[21]), .CO(
        dp_cluster_0_sub_487_C412_carry[22]), .S(s1_7_tmp_r[9]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_20 ( .A(dp_cluster_0_N77), .B(n1279), 
        .CI(dp_cluster_0_sub_487_C412_carry[20]), .CO(
        dp_cluster_0_sub_487_C412_carry[21]), .S(s1_7_tmp_r[8]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_19 ( .A(dp_cluster_0_N76), .B(n1280), 
        .CI(dp_cluster_0_sub_487_C412_carry[19]), .CO(
        dp_cluster_0_sub_487_C412_carry[20]), .S(s1_7_tmp_r[7]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_18 ( .A(dp_cluster_0_N75), .B(n1281), 
        .CI(dp_cluster_0_sub_487_C412_carry[18]), .CO(
        dp_cluster_0_sub_487_C412_carry[19]), .S(s1_7_tmp_r[6]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_17 ( .A(dp_cluster_0_N74), .B(n1282), 
        .CI(dp_cluster_0_sub_487_C412_carry[17]), .CO(
        dp_cluster_0_sub_487_C412_carry[18]), .S(s1_7_tmp_r[5]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_16 ( .A(dp_cluster_0_N73), .B(n1283), 
        .CI(dp_cluster_0_sub_487_C412_carry[16]), .CO(
        dp_cluster_0_sub_487_C412_carry[17]), .S(s1_7_tmp_r[4]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_15 ( .A(dp_cluster_2_N16), .B(n1251), 
        .CI(dp_cluster_2_sub_487_C409_carry[15]), .CO(
        dp_cluster_2_sub_487_C409_carry[16]), .S(s1_5_tmp_r[3]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_14 ( .A(dp_cluster_2_N15), .B(n1253), 
        .CI(dp_cluster_2_sub_487_C409_carry[14]), .CO(
        dp_cluster_2_sub_487_C409_carry[15]), .S(s1_5_tmp_r[2]) );
  FA1D0 dp_cluster_2_sub_487_C409_U2_13 ( .A(dp_cluster_2_N14), .B(n1254), 
        .CI(dp_cluster_2_sub_487_C409_carry[13]), .CO(
        dp_cluster_2_sub_487_C409_carry[14]), .S(s1_5_tmp_r[1]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_25 ( .A(dp_cluster_3_N138), .B(
        dp_cluster_3_N166), .CI(dp_cluster_3_add_514_C415_carry[25]), .CO(
        dp_cluster_3_add_514_C415_carry[26]), .S(s1_5_tmp_i[13]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_24 ( .A(dp_cluster_3_N137), .B(
        dp_cluster_3_N165), .CI(dp_cluster_3_add_514_C415_carry[24]), .CO(
        dp_cluster_3_add_514_C415_carry[25]), .S(s1_5_tmp_i[12]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_23 ( .A(dp_cluster_3_N136), .B(
        dp_cluster_3_N164), .CI(dp_cluster_3_add_514_C415_carry[23]), .CO(
        dp_cluster_3_add_514_C415_carry[24]), .S(s1_5_tmp_i[11]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_22 ( .A(dp_cluster_3_N135), .B(
        dp_cluster_3_N163), .CI(dp_cluster_3_add_514_C415_carry[22]), .CO(
        dp_cluster_3_add_514_C415_carry[23]), .S(s1_5_tmp_i[10]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_21 ( .A(dp_cluster_3_N134), .B(
        dp_cluster_3_N162), .CI(dp_cluster_3_add_514_C415_carry[21]), .CO(
        dp_cluster_3_add_514_C415_carry[22]), .S(s1_5_tmp_i[9]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_20 ( .A(dp_cluster_3_N133), .B(
        dp_cluster_3_N161), .CI(dp_cluster_3_add_514_C415_carry[20]), .CO(
        dp_cluster_3_add_514_C415_carry[21]), .S(s1_5_tmp_i[8]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_19 ( .A(dp_cluster_3_N132), .B(
        dp_cluster_3_N160), .CI(dp_cluster_3_add_514_C415_carry[19]), .CO(
        dp_cluster_3_add_514_C415_carry[20]), .S(s1_5_tmp_i[7]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_18 ( .A(dp_cluster_3_N131), .B(
        dp_cluster_3_N159), .CI(dp_cluster_3_add_514_C415_carry[18]), .CO(
        dp_cluster_3_add_514_C415_carry[19]), .S(s1_5_tmp_i[6]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_17 ( .A(dp_cluster_3_N130), .B(
        dp_cluster_3_N158), .CI(dp_cluster_3_add_514_C415_carry[17]), .CO(
        dp_cluster_3_add_514_C415_carry[18]), .S(s1_5_tmp_i[5]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_16 ( .A(dp_cluster_3_N129), .B(
        dp_cluster_3_N157), .CI(dp_cluster_3_add_514_C415_carry[16]), .CO(
        dp_cluster_3_add_514_C415_carry[17]), .S(s1_5_tmp_i[4]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_15 ( .A(dp_cluster_3_N128), .B(
        dp_cluster_3_N156), .CI(dp_cluster_3_add_514_C415_carry[15]), .CO(
        dp_cluster_3_add_514_C415_carry[16]), .S(s1_5_tmp_i[3]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_14 ( .A(dp_cluster_3_N127), .B(
        dp_cluster_3_N155), .CI(dp_cluster_3_add_514_C415_carry[14]), .CO(
        dp_cluster_3_add_514_C415_carry[15]), .S(s1_5_tmp_i[2]) );
  FA1D0 dp_cluster_3_add_514_C415_U1_13 ( .A(dp_cluster_3_N126), .B(
        dp_cluster_3_N154), .CI(dp_cluster_3_add_514_C415_carry[13]), .CO(
        dp_cluster_3_add_514_C415_carry[14]), .S(s1_5_tmp_i[1]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_15 ( .A(dp_cluster_0_N72), .B(n1284), 
        .CI(dp_cluster_0_sub_487_C412_carry[15]), .CO(
        dp_cluster_0_sub_487_C412_carry[16]), .S(s1_7_tmp_r[3]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_14 ( .A(dp_cluster_0_N71), .B(n1286), 
        .CI(dp_cluster_0_sub_487_C412_carry[14]), .CO(
        dp_cluster_0_sub_487_C412_carry[15]), .S(s1_7_tmp_r[2]) );
  FA1D0 dp_cluster_0_sub_487_C412_U2_13 ( .A(dp_cluster_0_N70), .B(n1287), 
        .CI(dp_cluster_0_sub_487_C412_carry[13]), .CO(
        dp_cluster_0_sub_487_C412_carry[14]), .S(s1_7_tmp_r[1]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_25 ( .A(dp_cluster_1_N194), .B(
        dp_cluster_1_N222), .CI(dp_cluster_1_add_514_C418_carry[25]), .CO(
        dp_cluster_1_add_514_C418_carry[26]), .S(s1_7_tmp_i[13]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_24 ( .A(dp_cluster_1_N193), .B(
        dp_cluster_1_N221), .CI(dp_cluster_1_add_514_C418_carry[24]), .CO(
        dp_cluster_1_add_514_C418_carry[25]), .S(s1_7_tmp_i[12]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_23 ( .A(dp_cluster_1_N192), .B(
        dp_cluster_1_N220), .CI(dp_cluster_1_add_514_C418_carry[23]), .CO(
        dp_cluster_1_add_514_C418_carry[24]), .S(s1_7_tmp_i[11]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_22 ( .A(dp_cluster_1_N191), .B(
        dp_cluster_1_N219), .CI(dp_cluster_1_add_514_C418_carry[22]), .CO(
        dp_cluster_1_add_514_C418_carry[23]), .S(s1_7_tmp_i[10]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_21 ( .A(dp_cluster_1_N190), .B(
        dp_cluster_1_N218), .CI(dp_cluster_1_add_514_C418_carry[21]), .CO(
        dp_cluster_1_add_514_C418_carry[22]), .S(s1_7_tmp_i[9]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_20 ( .A(dp_cluster_1_N189), .B(
        dp_cluster_1_N217), .CI(dp_cluster_1_add_514_C418_carry[20]), .CO(
        dp_cluster_1_add_514_C418_carry[21]), .S(s1_7_tmp_i[8]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_19 ( .A(dp_cluster_1_N188), .B(
        dp_cluster_1_N216), .CI(dp_cluster_1_add_514_C418_carry[19]), .CO(
        dp_cluster_1_add_514_C418_carry[20]), .S(s1_7_tmp_i[7]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_18 ( .A(dp_cluster_1_N187), .B(
        dp_cluster_1_N215), .CI(dp_cluster_1_add_514_C418_carry[18]), .CO(
        dp_cluster_1_add_514_C418_carry[19]), .S(s1_7_tmp_i[6]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_17 ( .A(dp_cluster_1_N186), .B(
        dp_cluster_1_N214), .CI(dp_cluster_1_add_514_C418_carry[17]), .CO(
        dp_cluster_1_add_514_C418_carry[18]), .S(s1_7_tmp_i[5]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_16 ( .A(dp_cluster_1_N185), .B(
        dp_cluster_1_N213), .CI(dp_cluster_1_add_514_C418_carry[16]), .CO(
        dp_cluster_1_add_514_C418_carry[17]), .S(s1_7_tmp_i[4]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_15 ( .A(dp_cluster_1_N184), .B(
        dp_cluster_1_N212), .CI(dp_cluster_1_add_514_C418_carry[15]), .CO(
        dp_cluster_1_add_514_C418_carry[16]), .S(s1_7_tmp_i[3]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_14 ( .A(dp_cluster_1_N183), .B(
        dp_cluster_1_N211), .CI(dp_cluster_1_add_514_C418_carry[14]), .CO(
        dp_cluster_1_add_514_C418_carry[15]), .S(s1_7_tmp_i[2]) );
  FA1D0 dp_cluster_1_add_514_C418_U1_13 ( .A(dp_cluster_1_N182), .B(
        dp_cluster_1_N210), .CI(dp_cluster_1_add_514_C418_carry[13]), .CO(
        dp_cluster_1_add_514_C418_carry[14]), .S(s1_7_tmp_i[1]) );
  TIEL U62 ( .ZN(xo7_i[1]) );
  TIEL U63 ( .ZN(xo7_i[2]) );
  TIEL U64 ( .ZN(xo7_i[3]) );
  TIEL U65 ( .ZN(xo7_i[4]) );
  TIEL U66 ( .ZN(xo7_i[5]) );
  TIEL U67 ( .ZN(xo7_i[6]) );
  TIEL U68 ( .ZN(xo7_i[7]) );
  TIEL U69 ( .ZN(xo7_i[8]) );
  TIEL U70 ( .ZN(xo7_i[9]) );
  TIEL U71 ( .ZN(xo7_i[10]) );
  TIEL U72 ( .ZN(xo7_i[11]) );
  TIEL U73 ( .ZN(xo7_i[12]) );
  TIEL U74 ( .ZN(xo7_i[13]) );
  TIEL U75 ( .ZN(xo7_i[14]) );
  TIEL U76 ( .ZN(xo7_i[15]) );
  TIEL U77 ( .ZN(xo7_i[16]) );
  TIEL U78 ( .ZN(xo7_i[17]) );
  TIEL U79 ( .ZN(xo7_i[18]) );
  TIEL U80 ( .ZN(xo7_i[19]) );
  TIEL U81 ( .ZN(xo7_i[20]) );
  TIEL U82 ( .ZN(xo7_i[21]) );
  TIEL U83 ( .ZN(xo7_i[22]) );
  TIEL U84 ( .ZN(xo7_i[23]) );
  TIEL U85 ( .ZN(xo7_i[24]) );
  TIEL U86 ( .ZN(xo7_i[25]) );
  TIEL U87 ( .ZN(xo7_i[26]) );
  TIEL U88 ( .ZN(xo7_i[27]) );
  TIEL U89 ( .ZN(xo7_i[28]) );
  TIEL U90 ( .ZN(xo7_i[29]) );
  TIEL U91 ( .ZN(xo7_i[30]) );
  TIEL U92 ( .ZN(xo7_i[31]) );
  TIEL U93 ( .ZN(xo7_i[32]) );
  TIEL U94 ( .ZN(xo7_i[33]) );
  TIEL U95 ( .ZN(xo7_i[34]) );
  TIEL U96 ( .ZN(xo7_i[35]) );
  TIEL U97 ( .ZN(xo7_i[36]) );
  TIEL U98 ( .ZN(xo7_i[37]) );
  TIEL U99 ( .ZN(xo7_i[38]) );
  TIEL U100 ( .ZN(xo7_i[39]) );
  TIEL U101 ( .ZN(xo7_i[40]) );
  TIEL U102 ( .ZN(xo7_i[41]) );
  TIEL U103 ( .ZN(xo7_i[42]) );
  TIEL U104 ( .ZN(xo7_i[43]) );
  TIEL U105 ( .ZN(xo7_i[44]) );
  TIEL U106 ( .ZN(xo7_i[45]) );
  TIEL U107 ( .ZN(xo7_i[46]) );
  TIEL U108 ( .ZN(xo7_i[47]) );
  TIEL U109 ( .ZN(xo6_i[0]) );
  TIEL U110 ( .ZN(xo6_i[1]) );
  TIEL U111 ( .ZN(xo6_i[2]) );
  TIEL U112 ( .ZN(xo6_i[3]) );
  TIEL U113 ( .ZN(xo6_i[4]) );
  TIEL U114 ( .ZN(xo6_i[5]) );
  TIEL U115 ( .ZN(xo6_i[6]) );
  TIEL U116 ( .ZN(xo6_i[7]) );
  TIEL U117 ( .ZN(xo6_i[8]) );
  TIEL U118 ( .ZN(xo6_i[9]) );
  TIEL U119 ( .ZN(xo6_i[10]) );
  TIEL U120 ( .ZN(xo6_i[11]) );
  TIEL U121 ( .ZN(xo6_i[12]) );
  TIEL U122 ( .ZN(xo6_i[13]) );
  TIEL U123 ( .ZN(xo6_i[14]) );
  TIEL U124 ( .ZN(xo6_i[15]) );
  TIEL U125 ( .ZN(xo6_i[16]) );
  TIEL U126 ( .ZN(xo6_i[17]) );
  TIEL U127 ( .ZN(xo6_i[18]) );
  TIEL U128 ( .ZN(xo6_i[19]) );
  TIEL U129 ( .ZN(xo6_i[20]) );
  TIEL U130 ( .ZN(xo6_i[21]) );
  TIEL U131 ( .ZN(xo6_i[22]) );
  TIEL U132 ( .ZN(xo6_i[23]) );
  TIEL U133 ( .ZN(xo6_i[24]) );
  TIEL U134 ( .ZN(xo6_i[25]) );
  TIEL U135 ( .ZN(xo6_i[26]) );
  TIEL U136 ( .ZN(xo6_i[27]) );
  TIEL U137 ( .ZN(xo6_i[28]) );
  TIEL U138 ( .ZN(xo6_i[29]) );
  TIEL U139 ( .ZN(xo6_i[30]) );
  TIEL U140 ( .ZN(xo6_i[31]) );
  TIEL U141 ( .ZN(xo6_i[32]) );
  TIEL U142 ( .ZN(xo6_i[33]) );
  TIEL U143 ( .ZN(xo6_i[34]) );
  TIEL U144 ( .ZN(xo6_i[35]) );
  TIEL U145 ( .ZN(xo6_i[36]) );
  TIEL U146 ( .ZN(xo6_i[37]) );
  TIEL U147 ( .ZN(xo6_i[38]) );
  TIEL U148 ( .ZN(xo6_i[39]) );
  TIEL U149 ( .ZN(xo6_i[40]) );
  TIEL U150 ( .ZN(xo6_i[41]) );
  TIEL U151 ( .ZN(xo6_i[42]) );
  TIEL U152 ( .ZN(xo6_i[43]) );
  TIEL U153 ( .ZN(xo6_i[44]) );
  TIEL U154 ( .ZN(xo6_i[45]) );
  TIEL U155 ( .ZN(xo6_i[46]) );
  TIEL U156 ( .ZN(xo6_i[47]) );
  TIEL U157 ( .ZN(xo5_i[0]) );
  TIEL U158 ( .ZN(xo5_i[1]) );
  TIEL U159 ( .ZN(xo5_i[2]) );
  TIEL U160 ( .ZN(xo5_i[3]) );
  TIEL U161 ( .ZN(xo5_i[4]) );
  TIEL U162 ( .ZN(xo5_i[5]) );
  TIEL U163 ( .ZN(xo5_i[6]) );
  TIEL U164 ( .ZN(xo5_i[7]) );
  TIEL U165 ( .ZN(xo5_i[8]) );
  TIEL U166 ( .ZN(xo5_i[9]) );
  TIEL U167 ( .ZN(xo5_i[10]) );
  TIEL U168 ( .ZN(xo5_i[11]) );
  TIEL U169 ( .ZN(xo5_i[12]) );
  TIEL U170 ( .ZN(xo5_i[13]) );
  TIEL U171 ( .ZN(xo5_i[14]) );
  TIEL U172 ( .ZN(xo5_i[15]) );
  TIEL U173 ( .ZN(xo5_i[16]) );
  TIEL U174 ( .ZN(xo5_i[17]) );
  TIEL U175 ( .ZN(xo5_i[18]) );
  TIEL U176 ( .ZN(xo5_i[19]) );
  TIEL U177 ( .ZN(xo5_i[20]) );
  TIEL U178 ( .ZN(xo5_i[21]) );
  TIEL U179 ( .ZN(xo5_i[22]) );
  TIEL U180 ( .ZN(xo5_i[23]) );
  TIEL U181 ( .ZN(xo5_i[24]) );
  TIEL U182 ( .ZN(xo5_i[25]) );
  TIEL U183 ( .ZN(xo5_i[26]) );
  TIEL U184 ( .ZN(xo5_i[27]) );
  TIEL U185 ( .ZN(xo5_i[28]) );
  TIEL U186 ( .ZN(xo5_i[29]) );
  TIEL U187 ( .ZN(xo5_i[30]) );
  TIEL U188 ( .ZN(xo5_i[31]) );
  TIEL U189 ( .ZN(xo5_i[32]) );
  TIEL U190 ( .ZN(xo5_i[33]) );
  TIEL U191 ( .ZN(xo5_i[34]) );
  TIEL U192 ( .ZN(xo5_i[35]) );
  TIEL U193 ( .ZN(xo5_i[36]) );
  TIEL U194 ( .ZN(xo5_i[37]) );
  TIEL U195 ( .ZN(xo5_i[38]) );
  TIEL U196 ( .ZN(xo5_i[39]) );
  TIEL U197 ( .ZN(xo5_i[40]) );
  TIEL U198 ( .ZN(xo5_i[41]) );
  TIEL U199 ( .ZN(xo5_i[42]) );
  TIEL U200 ( .ZN(xo5_i[43]) );
  TIEL U201 ( .ZN(xo5_i[44]) );
  TIEL U202 ( .ZN(xo5_i[45]) );
  TIEL U203 ( .ZN(xo5_i[46]) );
  TIEL U204 ( .ZN(xo5_i[47]) );
  TIEL U205 ( .ZN(xo4_i[0]) );
  TIEL U206 ( .ZN(xo4_i[1]) );
  TIEL U207 ( .ZN(xo4_i[2]) );
  TIEL U208 ( .ZN(xo4_i[3]) );
  TIEL U209 ( .ZN(xo4_i[4]) );
  TIEL U210 ( .ZN(xo4_i[5]) );
  TIEL U211 ( .ZN(xo4_i[6]) );
  TIEL U212 ( .ZN(xo4_i[7]) );
  TIEL U213 ( .ZN(xo4_i[8]) );
  TIEL U214 ( .ZN(xo4_i[9]) );
  TIEL U215 ( .ZN(xo4_i[10]) );
  TIEL U216 ( .ZN(xo4_i[11]) );
  TIEL U217 ( .ZN(xo4_i[12]) );
  TIEL U218 ( .ZN(xo4_i[13]) );
  TIEL U219 ( .ZN(xo4_i[14]) );
  TIEL U220 ( .ZN(xo4_i[15]) );
  TIEL U221 ( .ZN(xo4_i[16]) );
  TIEL U222 ( .ZN(xo4_i[17]) );
  TIEL U223 ( .ZN(xo4_i[18]) );
  TIEL U224 ( .ZN(xo4_i[19]) );
  TIEL U225 ( .ZN(xo4_i[20]) );
  TIEL U226 ( .ZN(xo4_i[21]) );
  TIEL U227 ( .ZN(xo4_i[22]) );
  TIEL U228 ( .ZN(xo4_i[23]) );
  TIEL U229 ( .ZN(xo4_i[24]) );
  TIEL U230 ( .ZN(xo4_i[25]) );
  TIEL U231 ( .ZN(xo4_i[26]) );
  TIEL U232 ( .ZN(xo4_i[27]) );
  TIEL U233 ( .ZN(xo4_i[28]) );
  TIEL U234 ( .ZN(xo4_i[29]) );
  TIEL U235 ( .ZN(xo4_i[30]) );
  TIEL U236 ( .ZN(xo4_i[31]) );
  TIEL U237 ( .ZN(xo4_i[32]) );
  TIEL U238 ( .ZN(xo4_i[33]) );
  TIEL U239 ( .ZN(xo4_i[34]) );
  TIEL U240 ( .ZN(xo4_i[35]) );
  TIEL U241 ( .ZN(xo4_i[36]) );
  TIEL U242 ( .ZN(xo4_i[37]) );
  TIEL U243 ( .ZN(xo4_i[38]) );
  TIEL U244 ( .ZN(xo4_i[39]) );
  TIEL U245 ( .ZN(xo4_i[40]) );
  TIEL U246 ( .ZN(xo4_i[41]) );
  TIEL U247 ( .ZN(xo4_i[42]) );
  TIEL U248 ( .ZN(xo4_i[43]) );
  TIEL U249 ( .ZN(xo4_i[44]) );
  TIEL U250 ( .ZN(xo4_i[45]) );
  TIEL U251 ( .ZN(xo4_i[46]) );
  TIEL U252 ( .ZN(xo4_i[47]) );
  TIEL U253 ( .ZN(xo3_i[0]) );
  TIEL U254 ( .ZN(xo3_i[1]) );
  TIEL U255 ( .ZN(xo3_i[2]) );
  TIEL U256 ( .ZN(xo3_i[3]) );
  TIEL U257 ( .ZN(xo3_i[4]) );
  TIEL U258 ( .ZN(xo3_i[5]) );
  TIEL U259 ( .ZN(xo3_i[6]) );
  TIEL U260 ( .ZN(xo3_i[7]) );
  TIEL U261 ( .ZN(xo3_i[8]) );
  TIEL U262 ( .ZN(xo3_i[9]) );
  TIEL U263 ( .ZN(xo3_i[10]) );
  TIEL U264 ( .ZN(xo3_i[11]) );
  TIEL U265 ( .ZN(xo3_i[12]) );
  TIEL U266 ( .ZN(xo3_i[13]) );
  TIEL U267 ( .ZN(xo3_i[14]) );
  TIEL U268 ( .ZN(xo3_i[15]) );
  TIEL U269 ( .ZN(xo3_i[16]) );
  TIEL U270 ( .ZN(xo3_i[17]) );
  TIEL U271 ( .ZN(xo3_i[18]) );
  TIEL U272 ( .ZN(xo3_i[19]) );
  TIEL U273 ( .ZN(xo3_i[20]) );
  TIEL U274 ( .ZN(xo3_i[21]) );
  TIEL U275 ( .ZN(xo3_i[22]) );
  TIEL U276 ( .ZN(xo3_i[23]) );
  TIEL U277 ( .ZN(xo3_i[24]) );
  TIEL U278 ( .ZN(xo3_i[25]) );
  TIEL U279 ( .ZN(xo3_i[26]) );
  TIEL U280 ( .ZN(xo3_i[27]) );
  TIEL U281 ( .ZN(xo3_i[28]) );
  TIEL U282 ( .ZN(xo3_i[29]) );
  TIEL U283 ( .ZN(xo3_i[30]) );
  TIEL U284 ( .ZN(xo3_i[31]) );
  TIEL U285 ( .ZN(xo3_i[32]) );
  TIEL U286 ( .ZN(xo3_i[33]) );
  TIEL U287 ( .ZN(xo3_i[34]) );
  TIEL U288 ( .ZN(xo3_i[35]) );
  TIEL U289 ( .ZN(xo3_i[36]) );
  TIEL U290 ( .ZN(xo3_i[37]) );
  TIEL U291 ( .ZN(xo3_i[38]) );
  TIEL U292 ( .ZN(xo3_i[39]) );
  TIEL U293 ( .ZN(xo3_i[40]) );
  TIEL U294 ( .ZN(xo3_i[41]) );
  TIEL U295 ( .ZN(xo3_i[42]) );
  TIEL U296 ( .ZN(xo3_i[43]) );
  TIEL U297 ( .ZN(xo3_i[44]) );
  TIEL U298 ( .ZN(xo3_i[45]) );
  TIEL U299 ( .ZN(xo3_i[46]) );
  TIEL U300 ( .ZN(xo3_i[47]) );
  TIEL U301 ( .ZN(xo2_i[0]) );
  TIEL U302 ( .ZN(xo2_i[1]) );
  TIEL U303 ( .ZN(xo2_i[2]) );
  TIEL U304 ( .ZN(xo2_i[3]) );
  TIEL U305 ( .ZN(xo2_i[4]) );
  TIEL U306 ( .ZN(xo2_i[5]) );
  TIEL U307 ( .ZN(xo2_i[6]) );
  TIEL U308 ( .ZN(xo2_i[7]) );
  TIEL U309 ( .ZN(xo2_i[8]) );
  TIEL U310 ( .ZN(xo2_i[9]) );
  TIEL U311 ( .ZN(xo2_i[10]) );
  TIEL U312 ( .ZN(xo2_i[11]) );
  TIEL U313 ( .ZN(xo2_i[12]) );
  TIEL U314 ( .ZN(xo2_i[13]) );
  TIEL U315 ( .ZN(xo2_i[14]) );
  TIEL U316 ( .ZN(xo2_i[15]) );
  TIEL U317 ( .ZN(xo2_i[16]) );
  TIEL U318 ( .ZN(xo2_i[17]) );
  TIEL U319 ( .ZN(xo2_i[18]) );
  TIEL U320 ( .ZN(xo2_i[19]) );
  TIEL U321 ( .ZN(xo2_i[20]) );
  TIEL U322 ( .ZN(xo2_i[21]) );
  TIEL U323 ( .ZN(xo2_i[22]) );
  TIEL U324 ( .ZN(xo2_i[23]) );
  TIEL U325 ( .ZN(xo2_i[24]) );
  TIEL U326 ( .ZN(xo2_i[25]) );
  TIEL U327 ( .ZN(xo2_i[26]) );
  TIEL U328 ( .ZN(xo2_i[27]) );
  TIEL U329 ( .ZN(xo2_i[28]) );
  TIEL U330 ( .ZN(xo2_i[29]) );
  TIEL U331 ( .ZN(xo2_i[30]) );
  TIEL U332 ( .ZN(xo2_i[31]) );
  TIEL U333 ( .ZN(xo2_i[32]) );
  TIEL U334 ( .ZN(xo2_i[33]) );
  TIEL U335 ( .ZN(xo2_i[34]) );
  TIEL U336 ( .ZN(xo2_i[35]) );
  TIEL U337 ( .ZN(xo2_i[36]) );
  TIEL U338 ( .ZN(xo2_i[37]) );
  TIEL U339 ( .ZN(xo2_i[38]) );
  TIEL U340 ( .ZN(xo2_i[39]) );
  TIEL U341 ( .ZN(xo2_i[40]) );
  TIEL U342 ( .ZN(xo2_i[41]) );
  TIEL U343 ( .ZN(xo2_i[42]) );
  TIEL U344 ( .ZN(xo2_i[43]) );
  TIEL U345 ( .ZN(xo2_i[44]) );
  TIEL U346 ( .ZN(xo2_i[45]) );
  TIEL U347 ( .ZN(xo2_i[46]) );
  TIEL U348 ( .ZN(xo2_i[47]) );
  TIEL U349 ( .ZN(xo1_i[0]) );
  TIEL U350 ( .ZN(xo1_i[1]) );
  TIEL U351 ( .ZN(xo1_i[2]) );
  TIEL U352 ( .ZN(xo1_i[3]) );
  TIEL U353 ( .ZN(xo1_i[4]) );
  TIEL U354 ( .ZN(xo1_i[5]) );
  TIEL U355 ( .ZN(xo1_i[6]) );
  TIEL U356 ( .ZN(xo1_i[7]) );
  TIEL U357 ( .ZN(xo1_i[8]) );
  TIEL U358 ( .ZN(xo1_i[9]) );
  TIEL U359 ( .ZN(xo1_i[10]) );
  TIEL U360 ( .ZN(xo1_i[11]) );
  TIEL U361 ( .ZN(xo1_i[12]) );
  TIEL U362 ( .ZN(xo1_i[13]) );
  TIEL U363 ( .ZN(xo1_i[14]) );
  TIEL U364 ( .ZN(xo1_i[15]) );
  TIEL U365 ( .ZN(xo1_i[16]) );
  TIEL U366 ( .ZN(xo1_i[17]) );
  TIEL U367 ( .ZN(xo1_i[18]) );
  TIEL U368 ( .ZN(xo1_i[19]) );
  TIEL U369 ( .ZN(xo1_i[20]) );
  TIEL U370 ( .ZN(xo1_i[21]) );
  TIEL U371 ( .ZN(xo1_i[22]) );
  TIEL U372 ( .ZN(xo1_i[23]) );
  TIEL U373 ( .ZN(xo1_i[24]) );
  TIEL U374 ( .ZN(xo1_i[25]) );
  TIEL U375 ( .ZN(xo1_i[26]) );
  TIEL U376 ( .ZN(xo1_i[27]) );
  TIEL U377 ( .ZN(xo1_i[28]) );
  TIEL U378 ( .ZN(xo1_i[29]) );
  TIEL U379 ( .ZN(xo1_i[30]) );
  TIEL U380 ( .ZN(xo1_i[31]) );
  TIEL U381 ( .ZN(xo1_i[32]) );
  TIEL U382 ( .ZN(xo1_i[33]) );
  TIEL U383 ( .ZN(xo1_i[34]) );
  TIEL U384 ( .ZN(xo1_i[35]) );
  TIEL U385 ( .ZN(xo1_i[36]) );
  TIEL U386 ( .ZN(xo1_i[37]) );
  TIEL U387 ( .ZN(xo1_i[38]) );
  TIEL U388 ( .ZN(xo1_i[39]) );
  TIEL U389 ( .ZN(xo1_i[40]) );
  TIEL U390 ( .ZN(xo1_i[41]) );
  TIEL U391 ( .ZN(xo1_i[42]) );
  TIEL U392 ( .ZN(xo1_i[43]) );
  TIEL U393 ( .ZN(xo1_i[44]) );
  TIEL U394 ( .ZN(xo1_i[45]) );
  TIEL U395 ( .ZN(xo1_i[46]) );
  TIEL U396 ( .ZN(xo1_i[47]) );
  TIEL U397 ( .ZN(xo0_i[0]) );
  TIEL U398 ( .ZN(xo0_i[1]) );
  TIEL U399 ( .ZN(xo0_i[2]) );
  TIEL U400 ( .ZN(xo0_i[3]) );
  TIEL U401 ( .ZN(xo0_i[4]) );
  TIEL U402 ( .ZN(xo0_i[5]) );
  TIEL U403 ( .ZN(xo0_i[6]) );
  TIEL U404 ( .ZN(xo0_i[7]) );
  TIEL U405 ( .ZN(xo0_i[8]) );
  TIEL U406 ( .ZN(xo0_i[9]) );
  TIEL U407 ( .ZN(xo0_i[10]) );
  TIEL U408 ( .ZN(xo0_i[11]) );
  TIEL U409 ( .ZN(xo0_i[12]) );
  TIEL U410 ( .ZN(xo0_i[13]) );
  TIEL U411 ( .ZN(xo0_i[14]) );
  TIEL U412 ( .ZN(xo0_i[15]) );
  TIEL U413 ( .ZN(xo0_i[16]) );
  TIEL U414 ( .ZN(xo0_i[17]) );
  TIEL U415 ( .ZN(xo0_i[18]) );
  TIEL U416 ( .ZN(xo0_i[19]) );
  TIEL U417 ( .ZN(xo0_i[20]) );
  TIEL U418 ( .ZN(xo0_i[21]) );
  TIEL U419 ( .ZN(xo0_i[22]) );
  TIEL U420 ( .ZN(xo0_i[23]) );
  TIEL U421 ( .ZN(xo0_i[24]) );
  TIEL U422 ( .ZN(xo0_i[25]) );
  TIEL U423 ( .ZN(xo0_i[26]) );
  TIEL U424 ( .ZN(xo0_i[27]) );
  TIEL U425 ( .ZN(xo0_i[28]) );
  TIEL U426 ( .ZN(xo0_i[29]) );
  TIEL U427 ( .ZN(xo0_i[30]) );
  TIEL U428 ( .ZN(xo0_i[31]) );
  TIEL U429 ( .ZN(xo0_i[32]) );
  TIEL U430 ( .ZN(xo0_i[33]) );
  TIEL U431 ( .ZN(xo0_i[34]) );
  TIEL U432 ( .ZN(xo0_i[35]) );
  TIEL U433 ( .ZN(xo0_i[36]) );
  TIEL U434 ( .ZN(xo0_i[37]) );
  TIEL U435 ( .ZN(xo0_i[38]) );
  TIEL U436 ( .ZN(xo0_i[39]) );
  TIEL U437 ( .ZN(xo0_i[40]) );
  TIEL U438 ( .ZN(xo0_i[41]) );
  TIEL U439 ( .ZN(xo0_i[42]) );
  TIEL U440 ( .ZN(xo0_i[43]) );
  TIEL U441 ( .ZN(xo0_i[44]) );
  TIEL U442 ( .ZN(xo0_i[45]) );
  TIEL U443 ( .ZN(xo0_i[46]) );
  TIEL U444 ( .ZN(xo0_i[47]) );
  TIEL U445 ( .ZN(xo7_r[0]) );
  TIEL U446 ( .ZN(xo7_r[1]) );
  TIEL U447 ( .ZN(xo7_r[2]) );
  TIEL U448 ( .ZN(xo7_r[3]) );
  TIEL U449 ( .ZN(xo7_r[4]) );
  TIEL U450 ( .ZN(xo7_r[5]) );
  TIEL U451 ( .ZN(xo7_r[6]) );
  TIEL U452 ( .ZN(xo7_r[7]) );
  TIEL U453 ( .ZN(xo7_r[8]) );
  TIEL U454 ( .ZN(xo7_r[9]) );
  TIEL U455 ( .ZN(xo7_r[10]) );
  TIEL U456 ( .ZN(xo7_r[11]) );
  TIEL U457 ( .ZN(xo7_r[12]) );
  TIEL U458 ( .ZN(xo7_r[13]) );
  TIEL U459 ( .ZN(xo7_r[14]) );
  TIEL U460 ( .ZN(xo7_r[15]) );
  TIEL U461 ( .ZN(xo7_r[16]) );
  TIEL U462 ( .ZN(xo7_r[17]) );
  TIEL U463 ( .ZN(xo7_r[18]) );
  TIEL U464 ( .ZN(xo7_r[19]) );
  TIEL U465 ( .ZN(xo7_r[20]) );
  TIEL U466 ( .ZN(xo7_r[21]) );
  TIEL U467 ( .ZN(xo7_r[22]) );
  TIEL U468 ( .ZN(xo7_r[23]) );
  TIEL U469 ( .ZN(xo7_r[24]) );
  TIEL U470 ( .ZN(xo7_r[25]) );
  TIEL U471 ( .ZN(xo7_r[26]) );
  TIEL U472 ( .ZN(xo7_r[27]) );
  TIEL U473 ( .ZN(xo7_r[28]) );
  TIEL U474 ( .ZN(xo7_r[29]) );
  TIEL U475 ( .ZN(xo7_r[30]) );
  TIEL U476 ( .ZN(xo7_r[31]) );
  TIEL U477 ( .ZN(xo7_r[32]) );
  TIEL U478 ( .ZN(xo7_r[33]) );
  TIEL U479 ( .ZN(xo7_r[34]) );
  TIEL U480 ( .ZN(xo7_r[35]) );
  TIEL U481 ( .ZN(xo7_r[36]) );
  TIEL U482 ( .ZN(xo7_r[37]) );
  TIEL U483 ( .ZN(xo7_r[38]) );
  TIEL U484 ( .ZN(xo7_r[39]) );
  TIEL U485 ( .ZN(xo7_r[40]) );
  TIEL U486 ( .ZN(xo7_r[41]) );
  TIEL U487 ( .ZN(xo7_r[42]) );
  TIEL U488 ( .ZN(xo7_r[43]) );
  TIEL U489 ( .ZN(xo7_r[44]) );
  TIEL U490 ( .ZN(xo7_r[45]) );
  TIEL U491 ( .ZN(xo7_r[46]) );
  TIEL U492 ( .ZN(xo7_r[47]) );
  TIEL U493 ( .ZN(xo6_r[0]) );
  TIEL U494 ( .ZN(xo6_r[1]) );
  TIEL U495 ( .ZN(xo6_r[2]) );
  TIEL U496 ( .ZN(xo6_r[3]) );
  TIEL U497 ( .ZN(xo6_r[4]) );
  TIEL U498 ( .ZN(xo6_r[5]) );
  TIEL U499 ( .ZN(xo6_r[6]) );
  TIEL U500 ( .ZN(xo6_r[7]) );
  TIEL U501 ( .ZN(xo6_r[8]) );
  TIEL U502 ( .ZN(xo6_r[9]) );
  TIEL U503 ( .ZN(xo6_r[10]) );
  TIEL U504 ( .ZN(xo6_r[11]) );
  TIEL U505 ( .ZN(xo6_r[12]) );
  TIEL U506 ( .ZN(xo6_r[13]) );
  TIEL U507 ( .ZN(xo6_r[14]) );
  TIEL U508 ( .ZN(xo6_r[15]) );
  TIEL U509 ( .ZN(xo6_r[16]) );
  TIEL U510 ( .ZN(xo6_r[17]) );
  TIEL U511 ( .ZN(xo6_r[18]) );
  TIEL U512 ( .ZN(xo6_r[19]) );
  TIEL U513 ( .ZN(xo6_r[20]) );
  TIEL U514 ( .ZN(xo6_r[21]) );
  TIEL U515 ( .ZN(xo6_r[22]) );
  TIEL U516 ( .ZN(xo6_r[23]) );
  TIEL U517 ( .ZN(xo6_r[24]) );
  TIEL U518 ( .ZN(xo6_r[25]) );
  TIEL U519 ( .ZN(xo6_r[26]) );
  TIEL U520 ( .ZN(xo6_r[27]) );
  TIEL U521 ( .ZN(xo6_r[28]) );
  TIEL U522 ( .ZN(xo6_r[29]) );
  TIEL U523 ( .ZN(xo6_r[30]) );
  TIEL U524 ( .ZN(xo6_r[31]) );
  TIEL U525 ( .ZN(xo6_r[32]) );
  TIEL U526 ( .ZN(xo6_r[33]) );
  TIEL U527 ( .ZN(xo6_r[34]) );
  TIEL U528 ( .ZN(xo6_r[35]) );
  TIEL U529 ( .ZN(xo6_r[36]) );
  TIEL U530 ( .ZN(xo6_r[37]) );
  TIEL U531 ( .ZN(xo6_r[38]) );
  TIEL U532 ( .ZN(xo6_r[39]) );
  TIEL U533 ( .ZN(xo6_r[40]) );
  TIEL U534 ( .ZN(xo6_r[41]) );
  TIEL U535 ( .ZN(xo6_r[42]) );
  TIEL U536 ( .ZN(xo6_r[43]) );
  TIEL U537 ( .ZN(xo6_r[44]) );
  TIEL U538 ( .ZN(xo6_r[45]) );
  TIEL U539 ( .ZN(xo6_r[46]) );
  TIEL U540 ( .ZN(xo6_r[47]) );
  TIEL U541 ( .ZN(xo5_r[0]) );
  TIEL U542 ( .ZN(xo5_r[1]) );
  TIEL U543 ( .ZN(xo5_r[2]) );
  TIEL U544 ( .ZN(xo5_r[3]) );
  TIEL U545 ( .ZN(xo5_r[4]) );
  TIEL U546 ( .ZN(xo5_r[5]) );
  TIEL U547 ( .ZN(xo5_r[6]) );
  TIEL U548 ( .ZN(xo5_r[7]) );
  TIEL U549 ( .ZN(xo5_r[8]) );
  TIEL U550 ( .ZN(xo5_r[9]) );
  TIEL U551 ( .ZN(xo5_r[10]) );
  TIEL U552 ( .ZN(xo5_r[11]) );
  TIEL U553 ( .ZN(xo5_r[12]) );
  TIEL U554 ( .ZN(xo5_r[13]) );
  TIEL U555 ( .ZN(xo5_r[14]) );
  TIEL U556 ( .ZN(xo5_r[15]) );
  TIEL U557 ( .ZN(xo5_r[16]) );
  TIEL U558 ( .ZN(xo5_r[17]) );
  TIEL U559 ( .ZN(xo5_r[18]) );
  TIEL U560 ( .ZN(xo5_r[19]) );
  TIEL U561 ( .ZN(xo5_r[20]) );
  TIEL U562 ( .ZN(xo5_r[21]) );
  TIEL U563 ( .ZN(xo5_r[22]) );
  TIEL U564 ( .ZN(xo5_r[23]) );
  TIEL U565 ( .ZN(xo5_r[24]) );
  TIEL U566 ( .ZN(xo5_r[25]) );
  TIEL U567 ( .ZN(xo5_r[26]) );
  TIEL U568 ( .ZN(xo5_r[27]) );
  TIEL U569 ( .ZN(xo5_r[28]) );
  TIEL U570 ( .ZN(xo5_r[29]) );
  TIEL U571 ( .ZN(xo5_r[30]) );
  TIEL U572 ( .ZN(xo5_r[31]) );
  TIEL U573 ( .ZN(xo5_r[32]) );
  TIEL U574 ( .ZN(xo5_r[33]) );
  TIEL U575 ( .ZN(xo5_r[34]) );
  TIEL U576 ( .ZN(xo5_r[35]) );
  TIEL U577 ( .ZN(xo5_r[36]) );
  TIEL U578 ( .ZN(xo5_r[37]) );
  TIEL U579 ( .ZN(xo5_r[38]) );
  TIEL U580 ( .ZN(xo5_r[39]) );
  TIEL U581 ( .ZN(xo5_r[40]) );
  TIEL U582 ( .ZN(xo5_r[41]) );
  TIEL U583 ( .ZN(xo5_r[42]) );
  TIEL U584 ( .ZN(xo5_r[43]) );
  TIEL U585 ( .ZN(xo5_r[44]) );
  TIEL U586 ( .ZN(xo5_r[45]) );
  TIEL U587 ( .ZN(xo5_r[46]) );
  TIEL U588 ( .ZN(xo5_r[47]) );
  TIEL U589 ( .ZN(xo4_r[0]) );
  TIEL U590 ( .ZN(xo4_r[1]) );
  TIEL U591 ( .ZN(xo4_r[2]) );
  TIEL U592 ( .ZN(xo4_r[3]) );
  TIEL U593 ( .ZN(xo4_r[4]) );
  TIEL U594 ( .ZN(xo4_r[5]) );
  TIEL U595 ( .ZN(xo4_r[6]) );
  TIEL U596 ( .ZN(xo4_r[7]) );
  TIEL U597 ( .ZN(xo4_r[8]) );
  TIEL U598 ( .ZN(xo4_r[9]) );
  TIEL U599 ( .ZN(xo4_r[10]) );
  TIEL U600 ( .ZN(xo4_r[11]) );
  TIEL U601 ( .ZN(xo4_r[12]) );
  TIEL U602 ( .ZN(xo4_r[13]) );
  TIEL U603 ( .ZN(xo4_r[14]) );
  TIEL U604 ( .ZN(xo4_r[15]) );
  TIEL U605 ( .ZN(xo4_r[16]) );
  TIEL U606 ( .ZN(xo4_r[17]) );
  TIEL U607 ( .ZN(xo4_r[18]) );
  TIEL U608 ( .ZN(xo4_r[19]) );
  TIEL U609 ( .ZN(xo4_r[20]) );
  TIEL U610 ( .ZN(xo4_r[21]) );
  TIEL U611 ( .ZN(xo4_r[22]) );
  TIEL U612 ( .ZN(xo4_r[23]) );
  TIEL U613 ( .ZN(xo4_r[24]) );
  TIEL U614 ( .ZN(xo4_r[25]) );
  TIEL U615 ( .ZN(xo4_r[26]) );
  TIEL U616 ( .ZN(xo4_r[27]) );
  TIEL U617 ( .ZN(xo4_r[28]) );
  TIEL U618 ( .ZN(xo4_r[29]) );
  TIEL U619 ( .ZN(xo4_r[30]) );
  TIEL U620 ( .ZN(xo4_r[31]) );
  TIEL U621 ( .ZN(xo4_r[32]) );
  TIEL U622 ( .ZN(xo4_r[33]) );
  TIEL U623 ( .ZN(xo4_r[34]) );
  TIEL U624 ( .ZN(xo4_r[35]) );
  TIEL U625 ( .ZN(xo4_r[36]) );
  TIEL U626 ( .ZN(xo4_r[37]) );
  TIEL U627 ( .ZN(xo4_r[38]) );
  TIEL U628 ( .ZN(xo4_r[39]) );
  TIEL U629 ( .ZN(xo4_r[40]) );
  TIEL U630 ( .ZN(xo4_r[41]) );
  TIEL U631 ( .ZN(xo4_r[42]) );
  TIEL U632 ( .ZN(xo4_r[43]) );
  TIEL U633 ( .ZN(xo4_r[44]) );
  TIEL U634 ( .ZN(xo4_r[45]) );
  TIEL U635 ( .ZN(xo4_r[46]) );
  TIEL U636 ( .ZN(xo4_r[47]) );
  TIEL U637 ( .ZN(xo3_r[0]) );
  TIEL U638 ( .ZN(xo3_r[1]) );
  TIEL U639 ( .ZN(xo3_r[2]) );
  TIEL U640 ( .ZN(xo3_r[3]) );
  TIEL U641 ( .ZN(xo3_r[4]) );
  TIEL U642 ( .ZN(xo3_r[5]) );
  TIEL U643 ( .ZN(xo3_r[6]) );
  TIEL U644 ( .ZN(xo3_r[7]) );
  TIEL U645 ( .ZN(xo3_r[8]) );
  TIEL U646 ( .ZN(xo3_r[9]) );
  TIEL U647 ( .ZN(xo3_r[10]) );
  TIEL U648 ( .ZN(xo3_r[11]) );
  TIEL U649 ( .ZN(xo3_r[12]) );
  TIEL U650 ( .ZN(xo3_r[13]) );
  TIEL U651 ( .ZN(xo3_r[14]) );
  TIEL U652 ( .ZN(xo3_r[15]) );
  TIEL U653 ( .ZN(xo3_r[16]) );
  TIEL U654 ( .ZN(xo3_r[17]) );
  TIEL U655 ( .ZN(xo3_r[18]) );
  TIEL U656 ( .ZN(xo3_r[19]) );
  TIEL U657 ( .ZN(xo3_r[20]) );
  TIEL U658 ( .ZN(xo3_r[21]) );
  TIEL U659 ( .ZN(xo3_r[22]) );
  TIEL U660 ( .ZN(xo3_r[23]) );
  TIEL U661 ( .ZN(xo3_r[24]) );
  TIEL U662 ( .ZN(xo3_r[25]) );
  TIEL U663 ( .ZN(xo3_r[26]) );
  TIEL U664 ( .ZN(xo3_r[27]) );
  TIEL U665 ( .ZN(xo3_r[28]) );
  TIEL U666 ( .ZN(xo3_r[29]) );
  TIEL U667 ( .ZN(xo3_r[30]) );
  TIEL U668 ( .ZN(xo3_r[31]) );
  TIEL U669 ( .ZN(xo3_r[32]) );
  TIEL U670 ( .ZN(xo3_r[33]) );
  TIEL U671 ( .ZN(xo3_r[34]) );
  TIEL U672 ( .ZN(xo3_r[35]) );
  TIEL U673 ( .ZN(xo3_r[36]) );
  TIEL U674 ( .ZN(xo3_r[37]) );
  TIEL U675 ( .ZN(xo3_r[38]) );
  TIEL U676 ( .ZN(xo3_r[39]) );
  TIEL U677 ( .ZN(xo3_r[40]) );
  TIEL U678 ( .ZN(xo3_r[41]) );
  TIEL U679 ( .ZN(xo3_r[42]) );
  TIEL U680 ( .ZN(xo3_r[43]) );
  TIEL U681 ( .ZN(xo3_r[44]) );
  TIEL U682 ( .ZN(xo3_r[45]) );
  TIEL U683 ( .ZN(xo3_r[46]) );
  TIEL U684 ( .ZN(xo3_r[47]) );
  TIEL U685 ( .ZN(xo2_r[0]) );
  TIEL U686 ( .ZN(xo2_r[1]) );
  TIEL U687 ( .ZN(xo2_r[2]) );
  TIEL U688 ( .ZN(xo2_r[3]) );
  TIEL U689 ( .ZN(xo2_r[4]) );
  TIEL U690 ( .ZN(xo2_r[5]) );
  TIEL U691 ( .ZN(xo2_r[6]) );
  TIEL U692 ( .ZN(xo2_r[7]) );
  TIEL U693 ( .ZN(xo2_r[8]) );
  TIEL U694 ( .ZN(xo2_r[9]) );
  TIEL U695 ( .ZN(xo2_r[10]) );
  TIEL U696 ( .ZN(xo2_r[11]) );
  TIEL U697 ( .ZN(xo2_r[12]) );
  TIEL U698 ( .ZN(xo2_r[13]) );
  TIEL U699 ( .ZN(xo2_r[14]) );
  TIEL U700 ( .ZN(xo2_r[15]) );
  TIEL U701 ( .ZN(xo2_r[16]) );
  TIEL U702 ( .ZN(xo2_r[17]) );
  TIEL U703 ( .ZN(xo2_r[18]) );
  TIEL U704 ( .ZN(xo2_r[19]) );
  TIEL U705 ( .ZN(xo2_r[20]) );
  TIEL U706 ( .ZN(xo2_r[21]) );
  TIEL U707 ( .ZN(xo2_r[22]) );
  TIEL U708 ( .ZN(xo2_r[23]) );
  TIEL U709 ( .ZN(xo2_r[24]) );
  TIEL U710 ( .ZN(xo2_r[25]) );
  TIEL U711 ( .ZN(xo2_r[26]) );
  TIEL U712 ( .ZN(xo2_r[27]) );
  TIEL U713 ( .ZN(xo2_r[28]) );
  TIEL U714 ( .ZN(xo2_r[29]) );
  TIEL U715 ( .ZN(xo2_r[30]) );
  TIEL U716 ( .ZN(xo2_r[31]) );
  TIEL U717 ( .ZN(xo2_r[32]) );
  TIEL U718 ( .ZN(xo2_r[33]) );
  TIEL U719 ( .ZN(xo2_r[34]) );
  TIEL U720 ( .ZN(xo2_r[35]) );
  TIEL U721 ( .ZN(xo2_r[36]) );
  TIEL U722 ( .ZN(xo2_r[37]) );
  TIEL U723 ( .ZN(xo2_r[38]) );
  TIEL U724 ( .ZN(xo2_r[39]) );
  TIEL U725 ( .ZN(xo2_r[40]) );
  TIEL U726 ( .ZN(xo2_r[41]) );
  TIEL U727 ( .ZN(xo2_r[42]) );
  TIEL U728 ( .ZN(xo2_r[43]) );
  TIEL U729 ( .ZN(xo2_r[44]) );
  TIEL U730 ( .ZN(xo2_r[45]) );
  TIEL U731 ( .ZN(xo2_r[46]) );
  TIEL U732 ( .ZN(xo2_r[47]) );
  TIEL U733 ( .ZN(xo1_r[0]) );
  TIEL U734 ( .ZN(xo1_r[1]) );
  TIEL U735 ( .ZN(xo1_r[2]) );
  TIEL U736 ( .ZN(xo1_r[3]) );
  TIEL U737 ( .ZN(xo1_r[4]) );
  TIEL U738 ( .ZN(xo1_r[5]) );
  TIEL U739 ( .ZN(xo1_r[6]) );
  TIEL U740 ( .ZN(xo1_r[7]) );
  TIEL U741 ( .ZN(xo1_r[8]) );
  TIEL U742 ( .ZN(xo1_r[9]) );
  TIEL U743 ( .ZN(xo1_r[10]) );
  TIEL U744 ( .ZN(xo1_r[11]) );
  TIEL U745 ( .ZN(xo1_r[12]) );
  TIEL U746 ( .ZN(xo1_r[13]) );
  TIEL U747 ( .ZN(xo1_r[14]) );
  TIEL U748 ( .ZN(xo1_r[15]) );
  TIEL U749 ( .ZN(xo1_r[16]) );
  TIEL U750 ( .ZN(xo1_r[17]) );
  TIEL U751 ( .ZN(xo1_r[18]) );
  TIEL U752 ( .ZN(xo1_r[19]) );
  TIEL U753 ( .ZN(xo1_r[20]) );
  TIEL U754 ( .ZN(xo1_r[21]) );
  TIEL U755 ( .ZN(xo1_r[22]) );
  TIEL U756 ( .ZN(xo1_r[23]) );
  TIEL U757 ( .ZN(xo1_r[24]) );
  TIEL U758 ( .ZN(xo1_r[25]) );
  TIEL U759 ( .ZN(xo1_r[26]) );
  TIEL U760 ( .ZN(xo1_r[27]) );
  TIEL U761 ( .ZN(xo1_r[28]) );
  TIEL U762 ( .ZN(xo1_r[29]) );
  TIEL U763 ( .ZN(xo1_r[30]) );
  TIEL U764 ( .ZN(xo1_r[31]) );
  TIEL U765 ( .ZN(xo1_r[32]) );
  TIEL U766 ( .ZN(xo1_r[33]) );
  TIEL U767 ( .ZN(xo1_r[34]) );
  TIEL U768 ( .ZN(xo1_r[35]) );
  TIEL U769 ( .ZN(xo1_r[36]) );
  TIEL U770 ( .ZN(xo1_r[37]) );
  TIEL U771 ( .ZN(xo1_r[38]) );
  TIEL U772 ( .ZN(xo1_r[39]) );
  TIEL U773 ( .ZN(xo1_r[40]) );
  TIEL U774 ( .ZN(xo1_r[41]) );
  TIEL U775 ( .ZN(xo1_r[42]) );
  TIEL U776 ( .ZN(xo1_r[43]) );
  TIEL U777 ( .ZN(xo1_r[44]) );
  TIEL U778 ( .ZN(xo1_r[45]) );
  TIEL U779 ( .ZN(xo1_r[46]) );
  TIEL U780 ( .ZN(xo1_r[47]) );
  TIEL U781 ( .ZN(xo0_r[0]) );
  TIEL U782 ( .ZN(xo0_r[1]) );
  TIEL U783 ( .ZN(xo0_r[2]) );
  TIEL U784 ( .ZN(xo0_r[3]) );
  TIEL U785 ( .ZN(xo0_r[4]) );
  TIEL U786 ( .ZN(xo0_r[5]) );
  TIEL U787 ( .ZN(xo0_r[6]) );
  TIEL U788 ( .ZN(xo0_r[7]) );
  TIEL U789 ( .ZN(xo0_r[8]) );
  TIEL U790 ( .ZN(xo0_r[9]) );
  TIEL U791 ( .ZN(xo0_r[10]) );
  TIEL U792 ( .ZN(xo0_r[11]) );
  TIEL U793 ( .ZN(xo0_r[12]) );
  TIEL U794 ( .ZN(xo0_r[13]) );
  TIEL U795 ( .ZN(xo0_r[14]) );
  TIEL U796 ( .ZN(xo0_r[15]) );
  TIEL U797 ( .ZN(xo0_r[16]) );
  TIEL U798 ( .ZN(xo0_r[17]) );
  TIEL U799 ( .ZN(xo0_r[18]) );
  TIEL U800 ( .ZN(xo0_r[19]) );
  TIEL U801 ( .ZN(xo0_r[20]) );
  TIEL U802 ( .ZN(xo0_r[21]) );
  TIEL U803 ( .ZN(xo0_r[22]) );
  TIEL U804 ( .ZN(xo0_r[23]) );
  TIEL U805 ( .ZN(xo0_r[24]) );
  TIEL U806 ( .ZN(xo0_r[25]) );
  TIEL U807 ( .ZN(xo0_r[26]) );
  TIEL U808 ( .ZN(xo0_r[27]) );
  TIEL U809 ( .ZN(xo0_r[28]) );
  TIEL U810 ( .ZN(xo0_r[29]) );
  TIEL U811 ( .ZN(xo0_r[30]) );
  TIEL U812 ( .ZN(xo0_r[31]) );
  TIEL U813 ( .ZN(xo0_r[32]) );
  TIEL U814 ( .ZN(xo0_r[33]) );
  TIEL U815 ( .ZN(xo0_r[34]) );
  TIEL U816 ( .ZN(xo0_r[35]) );
  TIEL U817 ( .ZN(xo0_r[36]) );
  TIEL U818 ( .ZN(xo0_r[37]) );
  TIEL U819 ( .ZN(xo0_r[38]) );
  TIEL U820 ( .ZN(xo0_r[39]) );
  TIEL U821 ( .ZN(xo0_r[40]) );
  TIEL U822 ( .ZN(xo0_r[41]) );
  TIEL U823 ( .ZN(xo0_r[42]) );
  TIEL U824 ( .ZN(xo0_r[43]) );
  TIEL U825 ( .ZN(xo0_r[44]) );
  TIEL U826 ( .ZN(xo0_r[45]) );
  TIEL U827 ( .ZN(xo0_r[46]) );
  TIEL U828 ( .ZN(xo0_r[47]) );
  XNR3D1 U829 ( .A1(n1837), .A2(n1836), .A3(n1835), .ZN(n905) );
  XNR3D1 U830 ( .A1(n2488), .A2(n2487), .A3(n2486), .ZN(n906) );
  AN2XD1 U831 ( .A1(s2_4_i[0]), .A2(s2_5_i[0]), .Z(n907) );
  AN2XD1 U832 ( .A1(s2_4_r[0]), .A2(s2_5_r[0]), .Z(n908) );
  AN2XD1 U833 ( .A1(s2_0_i[0]), .A2(s2_1_i[0]), .Z(n909) );
  AN2XD1 U834 ( .A1(s2_0_r[0]), .A2(s2_1_r[0]), .Z(n910) );
  AN2XD1 U835 ( .A1(s2_6_i[0]), .A2(s2_7_tmp_i_0_), .Z(n911) );
  AN2XD1 U836 ( .A1(s2_6_r[0]), .A2(s2_7_i[0]), .Z(n912) );
  AN2XD1 U837 ( .A1(s2_2_i[0]), .A2(s2_3_tmp_i_0_), .Z(n913) );
  AN2XD1 U838 ( .A1(s2_2_r[0]), .A2(s2_3_i[0]), .Z(n914) );
  AN2XD1 U839 ( .A1(xo4_i_w_d1r[0]), .A2(xo6_i_w_d1r[0]), .Z(n915) );
  AN2XD1 U840 ( .A1(xo4_r_w_d1r[0]), .A2(xo6_r_w_d1r[0]), .Z(n916) );
  AN2XD1 U841 ( .A1(xo0_i_w_d1r[0]), .A2(xo2_i_w_d1r[0]), .Z(n917) );
  AN2XD1 U842 ( .A1(xo0_r_w_d1r[0]), .A2(xo2_r_w_d1r[0]), .Z(n918) );
  AN2XD1 U843 ( .A1(xo5_i_w_d1r[0]), .A2(xo7_i_w_d1r[0]), .Z(n919) );
  AN2XD1 U844 ( .A1(xo1_i_w_d1r[0]), .A2(xo3_i_w_d1r[0]), .Z(n920) );
  AN2XD1 U845 ( .A1(xo5_r_w_d1r[0]), .A2(xo7_r_w_d1r[0]), .Z(n921) );
  AN2XD1 U846 ( .A1(xo1_r_w_d1r[0]), .A2(xo3_r_w_d1r[0]), .Z(n922) );
  INVD1 U847 ( .I(dp_cluster_0_N98), .ZN(n1287) );
  INVD1 U848 ( .I(dp_cluster_0_N99), .ZN(n1286) );
  INVD1 U849 ( .I(dp_cluster_0_N100), .ZN(n1284) );
  INVD1 U850 ( .I(dp_cluster_2_N42), .ZN(n1254) );
  INVD1 U851 ( .I(dp_cluster_2_N43), .ZN(n1253) );
  INVD1 U852 ( .I(dp_cluster_2_N44), .ZN(n1251) );
  INVD1 U853 ( .I(dp_cluster_0_N101), .ZN(n1283) );
  INVD1 U854 ( .I(dp_cluster_0_N102), .ZN(n1282) );
  INVD1 U855 ( .I(dp_cluster_0_N103), .ZN(n1281) );
  INVD1 U856 ( .I(dp_cluster_0_N104), .ZN(n1280) );
  INVD1 U857 ( .I(dp_cluster_0_N105), .ZN(n1279) );
  INVD1 U858 ( .I(dp_cluster_0_N106), .ZN(n1278) );
  INVD1 U859 ( .I(dp_cluster_0_N107), .ZN(n1277) );
  INVD1 U860 ( .I(dp_cluster_0_N108), .ZN(n1276) );
  INVD1 U861 ( .I(dp_cluster_0_N109), .ZN(n1275) );
  INVD1 U862 ( .I(dp_cluster_0_N110), .ZN(n1274) );
  INVD1 U863 ( .I(dp_cluster_2_N45), .ZN(n1250) );
  INVD1 U864 ( .I(dp_cluster_2_N46), .ZN(n1249) );
  INVD1 U865 ( .I(dp_cluster_2_N47), .ZN(n1248) );
  INVD1 U866 ( .I(dp_cluster_2_N48), .ZN(n1247) );
  INVD1 U867 ( .I(dp_cluster_2_N49), .ZN(n1246) );
  INVD1 U868 ( .I(dp_cluster_2_N50), .ZN(n1245) );
  INVD1 U869 ( .I(dp_cluster_2_N51), .ZN(n1244) );
  INVD1 U870 ( .I(dp_cluster_2_N52), .ZN(n1243) );
  INVD1 U871 ( .I(dp_cluster_2_N53), .ZN(n1242) );
  INVD1 U872 ( .I(dp_cluster_2_N54), .ZN(n1241) );
  NR2D1 U873 ( .A1(dp_cluster_0_N65), .A2(n2005), .ZN(n2004) );
  OAI22D1 U874 ( .A1(n2003), .A2(n1164), .B1(dp_cluster_0_N92), .B2(n2002), 
        .ZN(n2005) );
  NR2D1 U875 ( .A1(dp_cluster_2_N9), .A2(n2656), .ZN(n2655) );
  OAI22D1 U876 ( .A1(n2654), .A2(n1125), .B1(dp_cluster_2_N36), .B2(n2653), 
        .ZN(n2656) );
  NR2D1 U877 ( .A1(dp_cluster_0_N67), .A2(n2009), .ZN(n2008) );
  OAI22D1 U878 ( .A1(n2007), .A2(n1160), .B1(dp_cluster_0_N94), .B2(n2006), 
        .ZN(n2009) );
  NR2D1 U879 ( .A1(dp_cluster_2_N11), .A2(n2660), .ZN(n2659) );
  OAI22D1 U880 ( .A1(n2658), .A2(n1121), .B1(dp_cluster_2_N38), .B2(n2657), 
        .ZN(n2660) );
  OAI21D1 U881 ( .A1(dp_cluster_1_N179), .A2(n2334), .B(dp_cluster_1_N207), 
        .ZN(n2333) );
  OAI21D1 U882 ( .A1(dp_cluster_3_N123), .A2(n2985), .B(dp_cluster_3_N151), 
        .ZN(n2984) );
  FA1D0 U883 ( .A(dp_cluster_0_mult_486_C412_n175), .B(
        dp_cluster_0_mult_486_C412_n165), .CI(dp_cluster_0_mult_486_C412_n64), 
        .CO(dp_cluster_0_mult_486_C412_n63), .S(dp_cluster_0_N100) );
  FA1D0 U884 ( .A(dp_cluster_2_mult_486_C409_n175), .B(
        dp_cluster_2_mult_486_C409_n165), .CI(dp_cluster_2_mult_486_C409_n64), 
        .CO(dp_cluster_2_mult_486_C409_n63), .S(dp_cluster_2_N44) );
  FA1D0 U885 ( .A(dp_cluster_1_mult_512_C418_n175), .B(
        dp_cluster_1_mult_512_C418_n165), .CI(dp_cluster_1_mult_512_C418_n64), 
        .CO(dp_cluster_1_mult_512_C418_n63), .S(dp_cluster_1_N184) );
  FA1D0 U886 ( .A(dp_cluster_1_mult_513_C418_n175), .B(
        dp_cluster_1_mult_513_C418_n165), .CI(dp_cluster_1_mult_513_C418_n64), 
        .CO(dp_cluster_1_mult_513_C418_n63), .S(dp_cluster_1_N212) );
  FA1D0 U887 ( .A(dp_cluster_0_mult_486_C412_n164), .B(
        dp_cluster_0_mult_486_C412_n154), .CI(dp_cluster_0_mult_486_C412_n63), 
        .CO(dp_cluster_0_mult_486_C412_n62), .S(dp_cluster_0_N101) );
  FA1D0 U888 ( .A(dp_cluster_0_mult_485_C412_n175), .B(
        dp_cluster_0_mult_485_C412_n165), .CI(dp_cluster_0_mult_485_C412_n64), 
        .CO(dp_cluster_0_mult_485_C412_n63), .S(dp_cluster_0_N72) );
  FA1D0 U889 ( .A(dp_cluster_3_mult_512_C415_n175), .B(
        dp_cluster_3_mult_512_C415_n165), .CI(dp_cluster_3_mult_512_C415_n64), 
        .CO(dp_cluster_3_mult_512_C415_n63), .S(dp_cluster_3_N128) );
  FA1D0 U890 ( .A(dp_cluster_3_mult_513_C415_n175), .B(
        dp_cluster_3_mult_513_C415_n165), .CI(dp_cluster_3_mult_513_C415_n64), 
        .CO(dp_cluster_3_mult_513_C415_n63), .S(dp_cluster_3_N156) );
  FA1D0 U891 ( .A(dp_cluster_2_mult_486_C409_n164), .B(
        dp_cluster_2_mult_486_C409_n154), .CI(dp_cluster_2_mult_486_C409_n63), 
        .CO(dp_cluster_2_mult_486_C409_n62), .S(dp_cluster_2_N45) );
  FA1D0 U892 ( .A(dp_cluster_2_mult_485_C409_n175), .B(
        dp_cluster_2_mult_485_C409_n165), .CI(dp_cluster_2_mult_485_C409_n64), 
        .CO(dp_cluster_2_mult_485_C409_n63), .S(dp_cluster_2_N16) );
  FA1D0 U893 ( .A(dp_cluster_1_mult_512_C418_n164), .B(
        dp_cluster_1_mult_512_C418_n154), .CI(dp_cluster_1_mult_512_C418_n63), 
        .CO(dp_cluster_1_mult_512_C418_n62), .S(dp_cluster_1_N185) );
  FA1D0 U894 ( .A(dp_cluster_1_mult_513_C418_n164), .B(
        dp_cluster_1_mult_513_C418_n154), .CI(dp_cluster_1_mult_513_C418_n63), 
        .CO(dp_cluster_1_mult_513_C418_n62), .S(dp_cluster_1_N213) );
  FA1D0 U895 ( .A(dp_cluster_0_mult_486_C412_n153), .B(
        dp_cluster_0_mult_486_C412_n143), .CI(dp_cluster_0_mult_486_C412_n62), 
        .CO(dp_cluster_0_mult_486_C412_n61), .S(dp_cluster_0_N102) );
  FA1D0 U896 ( .A(dp_cluster_0_mult_485_C412_n164), .B(
        dp_cluster_0_mult_485_C412_n154), .CI(dp_cluster_0_mult_485_C412_n63), 
        .CO(dp_cluster_0_mult_485_C412_n62), .S(dp_cluster_0_N73) );
  FA1D0 U897 ( .A(dp_cluster_3_mult_512_C415_n164), .B(
        dp_cluster_3_mult_512_C415_n154), .CI(dp_cluster_3_mult_512_C415_n63), 
        .CO(dp_cluster_3_mult_512_C415_n62), .S(dp_cluster_3_N129) );
  FA1D0 U898 ( .A(dp_cluster_3_mult_513_C415_n164), .B(
        dp_cluster_3_mult_513_C415_n154), .CI(dp_cluster_3_mult_513_C415_n63), 
        .CO(dp_cluster_3_mult_513_C415_n62), .S(dp_cluster_3_N157) );
  FA1D0 U899 ( .A(dp_cluster_2_mult_486_C409_n153), .B(
        dp_cluster_2_mult_486_C409_n143), .CI(dp_cluster_2_mult_486_C409_n62), 
        .CO(dp_cluster_2_mult_486_C409_n61), .S(dp_cluster_2_N46) );
  FA1D0 U900 ( .A(dp_cluster_2_mult_485_C409_n164), .B(
        dp_cluster_2_mult_485_C409_n154), .CI(dp_cluster_2_mult_485_C409_n63), 
        .CO(dp_cluster_2_mult_485_C409_n62), .S(dp_cluster_2_N17) );
  FA1D0 U901 ( .A(dp_cluster_1_mult_512_C418_n153), .B(
        dp_cluster_1_mult_512_C418_n143), .CI(dp_cluster_1_mult_512_C418_n62), 
        .CO(dp_cluster_1_mult_512_C418_n61), .S(dp_cluster_1_N186) );
  FA1D0 U902 ( .A(dp_cluster_1_mult_513_C418_n153), .B(
        dp_cluster_1_mult_513_C418_n143), .CI(dp_cluster_1_mult_513_C418_n62), 
        .CO(dp_cluster_1_mult_513_C418_n61), .S(dp_cluster_1_N214) );
  FA1D0 U903 ( .A(dp_cluster_0_mult_486_C412_n142), .B(
        dp_cluster_0_mult_486_C412_n134), .CI(dp_cluster_0_mult_486_C412_n61), 
        .CO(dp_cluster_0_mult_486_C412_n60), .S(dp_cluster_0_N103) );
  FA1D0 U904 ( .A(dp_cluster_0_mult_485_C412_n153), .B(
        dp_cluster_0_mult_485_C412_n143), .CI(dp_cluster_0_mult_485_C412_n62), 
        .CO(dp_cluster_0_mult_485_C412_n61), .S(dp_cluster_0_N74) );
  FA1D0 U905 ( .A(dp_cluster_3_mult_512_C415_n153), .B(
        dp_cluster_3_mult_512_C415_n143), .CI(dp_cluster_3_mult_512_C415_n62), 
        .CO(dp_cluster_3_mult_512_C415_n61), .S(dp_cluster_3_N130) );
  FA1D0 U906 ( .A(dp_cluster_3_mult_513_C415_n153), .B(
        dp_cluster_3_mult_513_C415_n143), .CI(dp_cluster_3_mult_513_C415_n62), 
        .CO(dp_cluster_3_mult_513_C415_n61), .S(dp_cluster_3_N158) );
  FA1D0 U907 ( .A(dp_cluster_2_mult_486_C409_n142), .B(
        dp_cluster_2_mult_486_C409_n134), .CI(dp_cluster_2_mult_486_C409_n61), 
        .CO(dp_cluster_2_mult_486_C409_n60), .S(dp_cluster_2_N47) );
  FA1D0 U908 ( .A(dp_cluster_2_mult_485_C409_n153), .B(
        dp_cluster_2_mult_485_C409_n143), .CI(dp_cluster_2_mult_485_C409_n62), 
        .CO(dp_cluster_2_mult_485_C409_n61), .S(dp_cluster_2_N18) );
  FA1D0 U909 ( .A(dp_cluster_1_mult_512_C418_n142), .B(
        dp_cluster_1_mult_512_C418_n134), .CI(dp_cluster_1_mult_512_C418_n61), 
        .CO(dp_cluster_1_mult_512_C418_n60), .S(dp_cluster_1_N187) );
  FA1D0 U910 ( .A(dp_cluster_1_mult_513_C418_n142), .B(
        dp_cluster_1_mult_513_C418_n134), .CI(dp_cluster_1_mult_513_C418_n61), 
        .CO(dp_cluster_1_mult_513_C418_n60), .S(dp_cluster_1_N215) );
  FA1D0 U911 ( .A(dp_cluster_0_mult_486_C412_n133), .B(
        dp_cluster_0_mult_486_C412_n124), .CI(dp_cluster_0_mult_486_C412_n60), 
        .CO(dp_cluster_0_mult_486_C412_n59), .S(dp_cluster_0_N104) );
  FA1D0 U912 ( .A(dp_cluster_0_mult_485_C412_n142), .B(
        dp_cluster_0_mult_485_C412_n134), .CI(dp_cluster_0_mult_485_C412_n61), 
        .CO(dp_cluster_0_mult_485_C412_n60), .S(dp_cluster_0_N75) );
  FA1D0 U913 ( .A(dp_cluster_3_mult_512_C415_n142), .B(
        dp_cluster_3_mult_512_C415_n134), .CI(dp_cluster_3_mult_512_C415_n61), 
        .CO(dp_cluster_3_mult_512_C415_n60), .S(dp_cluster_3_N131) );
  FA1D0 U914 ( .A(dp_cluster_3_mult_513_C415_n142), .B(
        dp_cluster_3_mult_513_C415_n134), .CI(dp_cluster_3_mult_513_C415_n61), 
        .CO(dp_cluster_3_mult_513_C415_n60), .S(dp_cluster_3_N159) );
  FA1D0 U915 ( .A(dp_cluster_2_mult_486_C409_n133), .B(
        dp_cluster_2_mult_486_C409_n124), .CI(dp_cluster_2_mult_486_C409_n60), 
        .CO(dp_cluster_2_mult_486_C409_n59), .S(dp_cluster_2_N48) );
  FA1D0 U916 ( .A(dp_cluster_2_mult_485_C409_n142), .B(
        dp_cluster_2_mult_485_C409_n134), .CI(dp_cluster_2_mult_485_C409_n61), 
        .CO(dp_cluster_2_mult_485_C409_n60), .S(dp_cluster_2_N19) );
  FA1D0 U917 ( .A(dp_cluster_1_mult_512_C418_n133), .B(
        dp_cluster_1_mult_512_C418_n124), .CI(dp_cluster_1_mult_512_C418_n60), 
        .CO(dp_cluster_1_mult_512_C418_n59), .S(dp_cluster_1_N188) );
  FA1D0 U918 ( .A(dp_cluster_1_mult_513_C418_n133), .B(
        dp_cluster_1_mult_513_C418_n124), .CI(dp_cluster_1_mult_513_C418_n60), 
        .CO(dp_cluster_1_mult_513_C418_n59), .S(dp_cluster_1_N216) );
  FA1D0 U919 ( .A(dp_cluster_0_mult_486_C412_n123), .B(
        dp_cluster_0_mult_486_C412_n116), .CI(dp_cluster_0_mult_486_C412_n59), 
        .CO(dp_cluster_0_mult_486_C412_n58), .S(dp_cluster_0_N105) );
  FA1D0 U920 ( .A(dp_cluster_0_mult_485_C412_n133), .B(
        dp_cluster_0_mult_485_C412_n124), .CI(dp_cluster_0_mult_485_C412_n60), 
        .CO(dp_cluster_0_mult_485_C412_n59), .S(dp_cluster_0_N76) );
  FA1D0 U921 ( .A(dp_cluster_3_mult_512_C415_n133), .B(
        dp_cluster_3_mult_512_C415_n124), .CI(dp_cluster_3_mult_512_C415_n60), 
        .CO(dp_cluster_3_mult_512_C415_n59), .S(dp_cluster_3_N132) );
  FA1D0 U922 ( .A(dp_cluster_3_mult_513_C415_n133), .B(
        dp_cluster_3_mult_513_C415_n124), .CI(dp_cluster_3_mult_513_C415_n60), 
        .CO(dp_cluster_3_mult_513_C415_n59), .S(dp_cluster_3_N160) );
  FA1D0 U923 ( .A(dp_cluster_2_mult_486_C409_n123), .B(
        dp_cluster_2_mult_486_C409_n116), .CI(dp_cluster_2_mult_486_C409_n59), 
        .CO(dp_cluster_2_mult_486_C409_n58), .S(dp_cluster_2_N49) );
  FA1D0 U924 ( .A(dp_cluster_2_mult_485_C409_n133), .B(
        dp_cluster_2_mult_485_C409_n124), .CI(dp_cluster_2_mult_485_C409_n60), 
        .CO(dp_cluster_2_mult_485_C409_n59), .S(dp_cluster_2_N20) );
  FA1D0 U925 ( .A(dp_cluster_1_mult_512_C418_n123), .B(
        dp_cluster_1_mult_512_C418_n116), .CI(dp_cluster_1_mult_512_C418_n59), 
        .CO(dp_cluster_1_mult_512_C418_n58), .S(dp_cluster_1_N189) );
  FA1D0 U926 ( .A(dp_cluster_1_mult_513_C418_n123), .B(
        dp_cluster_1_mult_513_C418_n116), .CI(dp_cluster_1_mult_513_C418_n59), 
        .CO(dp_cluster_1_mult_513_C418_n58), .S(dp_cluster_1_N217) );
  FA1D0 U927 ( .A(dp_cluster_0_mult_486_C412_n115), .B(
        dp_cluster_0_mult_486_C412_n108), .CI(dp_cluster_0_mult_486_C412_n58), 
        .CO(dp_cluster_0_mult_486_C412_n57), .S(dp_cluster_0_N106) );
  FA1D0 U928 ( .A(dp_cluster_0_mult_485_C412_n123), .B(
        dp_cluster_0_mult_485_C412_n116), .CI(dp_cluster_0_mult_485_C412_n59), 
        .CO(dp_cluster_0_mult_485_C412_n58), .S(dp_cluster_0_N77) );
  FA1D0 U929 ( .A(dp_cluster_3_mult_512_C415_n123), .B(
        dp_cluster_3_mult_512_C415_n116), .CI(dp_cluster_3_mult_512_C415_n59), 
        .CO(dp_cluster_3_mult_512_C415_n58), .S(dp_cluster_3_N133) );
  FA1D0 U930 ( .A(dp_cluster_3_mult_513_C415_n123), .B(
        dp_cluster_3_mult_513_C415_n116), .CI(dp_cluster_3_mult_513_C415_n59), 
        .CO(dp_cluster_3_mult_513_C415_n58), .S(dp_cluster_3_N161) );
  FA1D0 U931 ( .A(dp_cluster_2_mult_486_C409_n115), .B(
        dp_cluster_2_mult_486_C409_n108), .CI(dp_cluster_2_mult_486_C409_n58), 
        .CO(dp_cluster_2_mult_486_C409_n57), .S(dp_cluster_2_N50) );
  FA1D0 U932 ( .A(dp_cluster_2_mult_485_C409_n123), .B(
        dp_cluster_2_mult_485_C409_n116), .CI(dp_cluster_2_mult_485_C409_n59), 
        .CO(dp_cluster_2_mult_485_C409_n58), .S(dp_cluster_2_N21) );
  FA1D0 U933 ( .A(dp_cluster_1_mult_512_C418_n115), .B(
        dp_cluster_1_mult_512_C418_n108), .CI(dp_cluster_1_mult_512_C418_n58), 
        .CO(dp_cluster_1_mult_512_C418_n57), .S(dp_cluster_1_N190) );
  FA1D0 U934 ( .A(dp_cluster_1_mult_513_C418_n115), .B(
        dp_cluster_1_mult_513_C418_n108), .CI(dp_cluster_1_mult_513_C418_n58), 
        .CO(dp_cluster_1_mult_513_C418_n57), .S(dp_cluster_1_N218) );
  FA1D0 U935 ( .A(dp_cluster_0_mult_486_C412_n107), .B(
        dp_cluster_0_mult_486_C412_n102), .CI(dp_cluster_0_mult_486_C412_n57), 
        .CO(dp_cluster_0_mult_486_C412_n56), .S(dp_cluster_0_N107) );
  FA1D0 U936 ( .A(dp_cluster_0_mult_485_C412_n115), .B(
        dp_cluster_0_mult_485_C412_n108), .CI(dp_cluster_0_mult_485_C412_n58), 
        .CO(dp_cluster_0_mult_485_C412_n57), .S(dp_cluster_0_N78) );
  FA1D0 U937 ( .A(dp_cluster_3_mult_512_C415_n115), .B(
        dp_cluster_3_mult_512_C415_n108), .CI(dp_cluster_3_mult_512_C415_n58), 
        .CO(dp_cluster_3_mult_512_C415_n57), .S(dp_cluster_3_N134) );
  FA1D0 U938 ( .A(dp_cluster_3_mult_513_C415_n115), .B(
        dp_cluster_3_mult_513_C415_n108), .CI(dp_cluster_3_mult_513_C415_n58), 
        .CO(dp_cluster_3_mult_513_C415_n57), .S(dp_cluster_3_N162) );
  FA1D0 U939 ( .A(dp_cluster_2_mult_486_C409_n107), .B(
        dp_cluster_2_mult_486_C409_n102), .CI(dp_cluster_2_mult_486_C409_n57), 
        .CO(dp_cluster_2_mult_486_C409_n56), .S(dp_cluster_2_N51) );
  FA1D0 U940 ( .A(dp_cluster_2_mult_485_C409_n115), .B(
        dp_cluster_2_mult_485_C409_n108), .CI(dp_cluster_2_mult_485_C409_n58), 
        .CO(dp_cluster_2_mult_485_C409_n57), .S(dp_cluster_2_N22) );
  FA1D0 U941 ( .A(dp_cluster_1_mult_512_C418_n107), .B(
        dp_cluster_1_mult_512_C418_n102), .CI(dp_cluster_1_mult_512_C418_n57), 
        .CO(dp_cluster_1_mult_512_C418_n56), .S(dp_cluster_1_N191) );
  FA1D0 U942 ( .A(dp_cluster_1_mult_513_C418_n107), .B(
        dp_cluster_1_mult_513_C418_n102), .CI(dp_cluster_1_mult_513_C418_n57), 
        .CO(dp_cluster_1_mult_513_C418_n56), .S(dp_cluster_1_N219) );
  FA1D0 U943 ( .A(dp_cluster_0_mult_486_C412_n101), .B(
        dp_cluster_0_mult_486_C412_n95), .CI(dp_cluster_0_mult_486_C412_n56), 
        .CO(dp_cluster_0_mult_486_C412_n55), .S(dp_cluster_0_N108) );
  FA1D0 U944 ( .A(dp_cluster_0_mult_485_C412_n107), .B(
        dp_cluster_0_mult_485_C412_n102), .CI(dp_cluster_0_mult_485_C412_n57), 
        .CO(dp_cluster_0_mult_485_C412_n56), .S(dp_cluster_0_N79) );
  FA1D0 U945 ( .A(dp_cluster_3_mult_512_C415_n107), .B(
        dp_cluster_3_mult_512_C415_n102), .CI(dp_cluster_3_mult_512_C415_n57), 
        .CO(dp_cluster_3_mult_512_C415_n56), .S(dp_cluster_3_N135) );
  FA1D0 U946 ( .A(dp_cluster_3_mult_513_C415_n107), .B(
        dp_cluster_3_mult_513_C415_n102), .CI(dp_cluster_3_mult_513_C415_n57), 
        .CO(dp_cluster_3_mult_513_C415_n56), .S(dp_cluster_3_N163) );
  FA1D0 U947 ( .A(dp_cluster_2_mult_486_C409_n101), .B(
        dp_cluster_2_mult_486_C409_n95), .CI(dp_cluster_2_mult_486_C409_n56), 
        .CO(dp_cluster_2_mult_486_C409_n55), .S(dp_cluster_2_N52) );
  FA1D0 U948 ( .A(dp_cluster_2_mult_485_C409_n107), .B(
        dp_cluster_2_mult_485_C409_n102), .CI(dp_cluster_2_mult_485_C409_n57), 
        .CO(dp_cluster_2_mult_485_C409_n56), .S(dp_cluster_2_N23) );
  FA1D0 U949 ( .A(dp_cluster_1_mult_512_C418_n101), .B(
        dp_cluster_1_mult_512_C418_n95), .CI(dp_cluster_1_mult_512_C418_n56), 
        .CO(dp_cluster_1_mult_512_C418_n55), .S(dp_cluster_1_N192) );
  FA1D0 U950 ( .A(dp_cluster_1_mult_513_C418_n101), .B(
        dp_cluster_1_mult_513_C418_n95), .CI(dp_cluster_1_mult_513_C418_n56), 
        .CO(dp_cluster_1_mult_513_C418_n55), .S(dp_cluster_1_N220) );
  FA1D0 U951 ( .A(dp_cluster_0_mult_486_C412_n94), .B(
        dp_cluster_0_mult_486_C412_n90), .CI(dp_cluster_0_mult_486_C412_n55), 
        .CO(dp_cluster_0_mult_486_C412_n54), .S(dp_cluster_0_N109) );
  FA1D0 U952 ( .A(dp_cluster_0_mult_485_C412_n101), .B(
        dp_cluster_0_mult_485_C412_n95), .CI(dp_cluster_0_mult_485_C412_n56), 
        .CO(dp_cluster_0_mult_485_C412_n55), .S(dp_cluster_0_N80) );
  FA1D0 U953 ( .A(dp_cluster_3_mult_512_C415_n101), .B(
        dp_cluster_3_mult_512_C415_n95), .CI(dp_cluster_3_mult_512_C415_n56), 
        .CO(dp_cluster_3_mult_512_C415_n55), .S(dp_cluster_3_N136) );
  FA1D0 U954 ( .A(dp_cluster_3_mult_513_C415_n101), .B(
        dp_cluster_3_mult_513_C415_n95), .CI(dp_cluster_3_mult_513_C415_n56), 
        .CO(dp_cluster_3_mult_513_C415_n55), .S(dp_cluster_3_N164) );
  FA1D0 U955 ( .A(dp_cluster_2_mult_486_C409_n94), .B(
        dp_cluster_2_mult_486_C409_n90), .CI(dp_cluster_2_mult_486_C409_n55), 
        .CO(dp_cluster_2_mult_486_C409_n54), .S(dp_cluster_2_N53) );
  FA1D0 U956 ( .A(dp_cluster_2_mult_485_C409_n101), .B(
        dp_cluster_2_mult_485_C409_n95), .CI(dp_cluster_2_mult_485_C409_n56), 
        .CO(dp_cluster_2_mult_485_C409_n55), .S(dp_cluster_2_N24) );
  FA1D0 U957 ( .A(dp_cluster_1_mult_512_C418_n94), .B(
        dp_cluster_1_mult_512_C418_n90), .CI(dp_cluster_1_mult_512_C418_n55), 
        .CO(dp_cluster_1_mult_512_C418_n54), .S(dp_cluster_1_N193) );
  FA1D0 U958 ( .A(dp_cluster_1_mult_513_C418_n94), .B(
        dp_cluster_1_mult_513_C418_n90), .CI(dp_cluster_1_mult_513_C418_n55), 
        .CO(dp_cluster_1_mult_513_C418_n54), .S(dp_cluster_1_N221) );
  FA1D0 U959 ( .A(dp_cluster_0_mult_486_C412_n89), .B(
        dp_cluster_0_mult_486_C412_n85), .CI(dp_cluster_0_mult_486_C412_n54), 
        .CO(dp_cluster_0_mult_486_C412_n53), .S(dp_cluster_0_N110) );
  FA1D0 U960 ( .A(dp_cluster_0_mult_485_C412_n94), .B(
        dp_cluster_0_mult_485_C412_n90), .CI(dp_cluster_0_mult_485_C412_n55), 
        .CO(dp_cluster_0_mult_485_C412_n54), .S(dp_cluster_0_N81) );
  FA1D0 U961 ( .A(dp_cluster_3_mult_512_C415_n94), .B(
        dp_cluster_3_mult_512_C415_n90), .CI(dp_cluster_3_mult_512_C415_n55), 
        .CO(dp_cluster_3_mult_512_C415_n54), .S(dp_cluster_3_N137) );
  FA1D0 U962 ( .A(dp_cluster_3_mult_513_C415_n94), .B(
        dp_cluster_3_mult_513_C415_n90), .CI(dp_cluster_3_mult_513_C415_n55), 
        .CO(dp_cluster_3_mult_513_C415_n54), .S(dp_cluster_3_N165) );
  FA1D0 U963 ( .A(dp_cluster_2_mult_486_C409_n89), .B(
        dp_cluster_2_mult_486_C409_n85), .CI(dp_cluster_2_mult_486_C409_n54), 
        .CO(dp_cluster_2_mult_486_C409_n53), .S(dp_cluster_2_N54) );
  FA1D0 U964 ( .A(dp_cluster_2_mult_485_C409_n94), .B(
        dp_cluster_2_mult_485_C409_n90), .CI(dp_cluster_2_mult_485_C409_n55), 
        .CO(dp_cluster_2_mult_485_C409_n54), .S(dp_cluster_2_N25) );
  FA1D0 U965 ( .A(dp_cluster_1_mult_512_C418_n89), .B(
        dp_cluster_1_mult_512_C418_n85), .CI(dp_cluster_1_mult_512_C418_n54), 
        .CO(dp_cluster_1_mult_512_C418_n53), .S(dp_cluster_1_N194) );
  FA1D0 U966 ( .A(dp_cluster_1_mult_513_C418_n89), .B(
        dp_cluster_1_mult_513_C418_n85), .CI(dp_cluster_1_mult_513_C418_n54), 
        .CO(dp_cluster_1_mult_513_C418_n53), .S(dp_cluster_1_N222) );
  FA1D0 U967 ( .A(dp_cluster_0_mult_485_C412_n89), .B(
        dp_cluster_0_mult_485_C412_n85), .CI(dp_cluster_0_mult_485_C412_n54), 
        .CO(dp_cluster_0_mult_485_C412_n53), .S(dp_cluster_0_N82) );
  FA1D0 U968 ( .A(dp_cluster_3_mult_512_C415_n89), .B(
        dp_cluster_3_mult_512_C415_n85), .CI(dp_cluster_3_mult_512_C415_n54), 
        .CO(dp_cluster_3_mult_512_C415_n53), .S(dp_cluster_3_N138) );
  FA1D0 U969 ( .A(dp_cluster_3_mult_513_C415_n89), .B(
        dp_cluster_3_mult_513_C415_n85), .CI(dp_cluster_3_mult_513_C415_n54), 
        .CO(dp_cluster_3_mult_513_C415_n53), .S(dp_cluster_3_N166) );
  FA1D0 U970 ( .A(dp_cluster_2_mult_485_C409_n89), .B(
        dp_cluster_2_mult_485_C409_n85), .CI(dp_cluster_2_mult_485_C409_n54), 
        .CO(dp_cluster_2_mult_485_C409_n53), .S(dp_cluster_2_N26) );
  IOA21D1 U971 ( .A1(n2336), .A2(dp_cluster_1_N180), .B(n2335), .ZN(
        dp_cluster_1_add_514_C418_carry[12]) );
  OAI21D1 U972 ( .A1(dp_cluster_1_N180), .A2(n2336), .B(dp_cluster_1_N208), 
        .ZN(n2335) );
  IOA21D1 U973 ( .A1(n2334), .A2(dp_cluster_1_N179), .B(n2333), .ZN(n2336) );
  OAI22D1 U974 ( .A1(n2011), .A2(n1155), .B1(dp_cluster_0_N96), .B2(n2010), 
        .ZN(dp_cluster_0_sub_487_C412_carry[12]) );
  INVD1 U975 ( .I(dp_cluster_0_N97), .ZN(n1289) );
  IOA21D1 U976 ( .A1(n2987), .A2(dp_cluster_3_N124), .B(n2986), .ZN(
        dp_cluster_3_add_514_C415_carry[12]) );
  OAI21D1 U977 ( .A1(dp_cluster_3_N124), .A2(n2987), .B(dp_cluster_3_N152), 
        .ZN(n2986) );
  IOA21D1 U978 ( .A1(n2985), .A2(dp_cluster_3_N123), .B(n2984), .ZN(n2987) );
  OAI22D1 U979 ( .A1(n2662), .A2(n1116), .B1(dp_cluster_2_N40), .B2(n2661), 
        .ZN(dp_cluster_2_sub_487_C409_carry[12]) );
  INVD1 U980 ( .I(dp_cluster_2_N41), .ZN(n1256) );
  FA1D0 U981 ( .A(dp_cluster_0_mult_486_C412_n185), .B(
        dp_cluster_0_mult_486_C412_n194), .CI(dp_cluster_0_mult_486_C412_n66), 
        .CO(dp_cluster_0_mult_486_C412_n65), .S(dp_cluster_0_N98) );
  FA1D0 U982 ( .A(dp_cluster_2_mult_486_C409_n185), .B(
        dp_cluster_2_mult_486_C409_n194), .CI(dp_cluster_2_mult_486_C409_n66), 
        .CO(dp_cluster_2_mult_486_C409_n65), .S(dp_cluster_2_N42) );
  FA1D0 U983 ( .A(dp_cluster_1_mult_512_C418_n185), .B(
        dp_cluster_1_mult_512_C418_n194), .CI(dp_cluster_1_mult_512_C418_n66), 
        .CO(dp_cluster_1_mult_512_C418_n65), .S(dp_cluster_1_N182) );
  FA1D0 U984 ( .A(dp_cluster_1_mult_513_C418_n185), .B(
        dp_cluster_1_mult_513_C418_n194), .CI(dp_cluster_1_mult_513_C418_n66), 
        .CO(dp_cluster_1_mult_513_C418_n65), .S(dp_cluster_1_N210) );
  FA1D0 U985 ( .A(dp_cluster_0_mult_486_C412_n176), .B(
        dp_cluster_0_mult_486_C412_n184), .CI(dp_cluster_0_mult_486_C412_n65), 
        .CO(dp_cluster_0_mult_486_C412_n64), .S(dp_cluster_0_N99) );
  FA1D0 U986 ( .A(dp_cluster_0_mult_485_C412_n185), .B(
        dp_cluster_0_mult_485_C412_n194), .CI(dp_cluster_0_mult_485_C412_n66), 
        .CO(dp_cluster_0_mult_485_C412_n65), .S(dp_cluster_0_N70) );
  FA1D0 U987 ( .A(dp_cluster_3_mult_512_C415_n185), .B(
        dp_cluster_3_mult_512_C415_n194), .CI(dp_cluster_3_mult_512_C415_n66), 
        .CO(dp_cluster_3_mult_512_C415_n65), .S(dp_cluster_3_N126) );
  FA1D0 U988 ( .A(dp_cluster_3_mult_513_C415_n185), .B(
        dp_cluster_3_mult_513_C415_n194), .CI(dp_cluster_3_mult_513_C415_n66), 
        .CO(dp_cluster_3_mult_513_C415_n65), .S(dp_cluster_3_N154) );
  FA1D0 U989 ( .A(dp_cluster_2_mult_486_C409_n176), .B(
        dp_cluster_2_mult_486_C409_n184), .CI(dp_cluster_2_mult_486_C409_n65), 
        .CO(dp_cluster_2_mult_486_C409_n64), .S(dp_cluster_2_N43) );
  FA1D0 U990 ( .A(dp_cluster_2_mult_485_C409_n185), .B(
        dp_cluster_2_mult_485_C409_n194), .CI(dp_cluster_2_mult_485_C409_n66), 
        .CO(dp_cluster_2_mult_485_C409_n65), .S(dp_cluster_2_N14) );
  FA1D0 U991 ( .A(dp_cluster_1_mult_512_C418_n176), .B(
        dp_cluster_1_mult_512_C418_n184), .CI(dp_cluster_1_mult_512_C418_n65), 
        .CO(dp_cluster_1_mult_512_C418_n64), .S(dp_cluster_1_N183) );
  FA1D0 U992 ( .A(dp_cluster_1_mult_513_C418_n176), .B(
        dp_cluster_1_mult_513_C418_n184), .CI(dp_cluster_1_mult_513_C418_n65), 
        .CO(dp_cluster_1_mult_513_C418_n64), .S(dp_cluster_1_N211) );
  FA1D0 U993 ( .A(dp_cluster_0_mult_485_C412_n176), .B(
        dp_cluster_0_mult_485_C412_n184), .CI(dp_cluster_0_mult_485_C412_n65), 
        .CO(dp_cluster_0_mult_485_C412_n64), .S(dp_cluster_0_N71) );
  FA1D0 U994 ( .A(dp_cluster_3_mult_512_C415_n176), .B(
        dp_cluster_3_mult_512_C415_n184), .CI(dp_cluster_3_mult_512_C415_n65), 
        .CO(dp_cluster_3_mult_512_C415_n64), .S(dp_cluster_3_N127) );
  FA1D0 U995 ( .A(dp_cluster_3_mult_513_C415_n176), .B(
        dp_cluster_3_mult_513_C415_n184), .CI(dp_cluster_3_mult_513_C415_n65), 
        .CO(dp_cluster_3_mult_513_C415_n64), .S(dp_cluster_3_N155) );
  FA1D0 U996 ( .A(dp_cluster_2_mult_485_C409_n176), .B(
        dp_cluster_2_mult_485_C409_n184), .CI(dp_cluster_2_mult_485_C409_n65), 
        .CO(dp_cluster_2_mult_485_C409_n64), .S(dp_cluster_2_N15) );
  IOA21D1 U997 ( .A1(n2328), .A2(dp_cluster_1_N176), .B(n2327), .ZN(n2330) );
  OAI21D1 U998 ( .A1(dp_cluster_1_N176), .A2(n2328), .B(dp_cluster_1_N204), 
        .ZN(n2327) );
  IOA21D1 U999 ( .A1(n2326), .A2(dp_cluster_1_N175), .B(n2325), .ZN(n2328) );
  OAI21D1 U1000 ( .A1(dp_cluster_1_N175), .A2(n2326), .B(dp_cluster_1_N203), 
        .ZN(n2325) );
  IOA21D1 U1001 ( .A1(n2979), .A2(dp_cluster_3_N120), .B(n2978), .ZN(n2981) );
  OAI21D1 U1002 ( .A1(dp_cluster_3_N120), .A2(n2979), .B(dp_cluster_3_N148), 
        .ZN(n2978) );
  IOA21D1 U1003 ( .A1(n2977), .A2(dp_cluster_3_N119), .B(n2976), .ZN(n2979) );
  OAI21D1 U1004 ( .A1(dp_cluster_3_N119), .A2(n2977), .B(dp_cluster_3_N147), 
        .ZN(n2976) );
  IOA21D1 U1005 ( .A1(n2332), .A2(dp_cluster_1_N178), .B(n2331), .ZN(n2334) );
  OAI21D1 U1006 ( .A1(dp_cluster_1_N178), .A2(n2332), .B(dp_cluster_1_N206), 
        .ZN(n2331) );
  IOA21D1 U1007 ( .A1(n2330), .A2(dp_cluster_1_N177), .B(n2329), .ZN(n2332) );
  OAI21D1 U1008 ( .A1(dp_cluster_1_N177), .A2(n2330), .B(dp_cluster_1_N205), 
        .ZN(n2329) );
  IOA21D1 U1009 ( .A1(n2983), .A2(dp_cluster_3_N122), .B(n2982), .ZN(n2985) );
  OAI21D1 U1010 ( .A1(dp_cluster_3_N122), .A2(n2983), .B(dp_cluster_3_N150), 
        .ZN(n2982) );
  IOA21D1 U1011 ( .A1(n2981), .A2(dp_cluster_3_N121), .B(n2980), .ZN(n2983) );
  OAI21D1 U1012 ( .A1(dp_cluster_3_N121), .A2(n2981), .B(dp_cluster_3_N149), 
        .ZN(n2980) );
  INVD1 U1013 ( .I(dp_cluster_0_N62), .ZN(n1167) );
  INVD1 U1014 ( .I(dp_cluster_2_N6), .ZN(n1128) );
  INVD1 U1015 ( .I(dp_cluster_0_N64), .ZN(n1164) );
  INVD1 U1016 ( .I(dp_cluster_2_N8), .ZN(n1125) );
  INVD1 U1017 ( .I(dp_cluster_0_N66), .ZN(n1160) );
  INVD1 U1018 ( .I(dp_cluster_2_N10), .ZN(n1121) );
  INVD1 U1019 ( .I(dp_cluster_0_N68), .ZN(n1155) );
  INVD1 U1020 ( .I(dp_cluster_2_N12), .ZN(n1116) );
  INVD1 U1021 ( .I(dp_cluster_0_N111), .ZN(n1273) );
  INVD1 U1022 ( .I(dp_cluster_2_N55), .ZN(n1240) );
  OAI22D1 U1023 ( .A1(n2202), .A2(n971), .B1(n2300), .B2(n2201), .ZN(
        dp_cluster_1_mult_512_C418_n112) );
  OAI22D1 U1024 ( .A1(n2050), .A2(n965), .B1(n2148), .B2(n2049), .ZN(
        dp_cluster_1_mult_513_C418_n112) );
  OAI22D1 U1025 ( .A1(n1724), .A2(n953), .B1(n1822), .B2(n1723), .ZN(
        dp_cluster_0_mult_486_C412_n112) );
  OAI22D1 U1026 ( .A1(n1876), .A2(n959), .B1(n1974), .B2(n1875), .ZN(
        dp_cluster_0_mult_485_C412_n112) );
  OAI22D1 U1027 ( .A1(n2853), .A2(n995), .B1(n2951), .B2(n2852), .ZN(
        dp_cluster_3_mult_512_C415_n112) );
  OAI22D1 U1028 ( .A1(n2701), .A2(n989), .B1(n2799), .B2(n2700), .ZN(
        dp_cluster_3_mult_513_C415_n112) );
  OAI22D1 U1029 ( .A1(n2375), .A2(n977), .B1(n2473), .B2(n2374), .ZN(
        dp_cluster_2_mult_486_C409_n112) );
  OAI22D1 U1030 ( .A1(n2527), .A2(n983), .B1(n2625), .B2(n2526), .ZN(
        dp_cluster_2_mult_485_C409_n112) );
  NR2D1 U1031 ( .A1(dp_cluster_0_N63), .A2(n2001), .ZN(n2000) );
  OAI22D1 U1032 ( .A1(n1999), .A2(n1167), .B1(dp_cluster_0_N90), .B2(n1998), 
        .ZN(n2001) );
  NR2D1 U1033 ( .A1(dp_cluster_2_N7), .A2(n2652), .ZN(n2651) );
  OAI22D1 U1034 ( .A1(n2650), .A2(n1128), .B1(dp_cluster_2_N34), .B2(n2649), 
        .ZN(n2652) );
  FA1D0 U1035 ( .A(dp_cluster_1_mult_513_C418_n325), .B(
        dp_cluster_1_mult_513_C418_n339), .CI(dp_cluster_1_mult_513_C418_n353), 
        .CO(dp_cluster_1_mult_513_C418_n218), .S(
        dp_cluster_1_mult_513_C418_n219) );
  OAI22D1 U1036 ( .A1(n2120), .A2(n967), .B1(n2128), .B2(n2119), .ZN(
        dp_cluster_1_mult_513_C418_n353) );
  OAI22D1 U1037 ( .A1(n2104), .A2(n966), .B1(n2110), .B2(n2103), .ZN(
        dp_cluster_1_mult_513_C418_n339) );
  OAI22D1 U1038 ( .A1(n2088), .A2(n968), .B1(n2092), .B2(n2087), .ZN(
        dp_cluster_1_mult_513_C418_n325) );
  FA1D0 U1039 ( .A(dp_cluster_3_mult_513_C415_n325), .B(
        dp_cluster_3_mult_513_C415_n339), .CI(dp_cluster_3_mult_513_C415_n353), 
        .CO(dp_cluster_3_mult_513_C415_n218), .S(
        dp_cluster_3_mult_513_C415_n219) );
  OAI22D1 U1040 ( .A1(n2771), .A2(n991), .B1(n2779), .B2(n2770), .ZN(
        dp_cluster_3_mult_513_C415_n353) );
  OAI22D1 U1041 ( .A1(n2755), .A2(n990), .B1(n2761), .B2(n2754), .ZN(
        dp_cluster_3_mult_513_C415_n339) );
  OAI22D1 U1042 ( .A1(n2739), .A2(n992), .B1(n2743), .B2(n2738), .ZN(
        dp_cluster_3_mult_513_C415_n325) );
  FA1D0 U1043 ( .A(dp_cluster_1_mult_512_C418_n325), .B(
        dp_cluster_1_mult_512_C418_n339), .CI(dp_cluster_1_mult_512_C418_n353), 
        .CO(dp_cluster_1_mult_512_C418_n218), .S(
        dp_cluster_1_mult_512_C418_n219) );
  OAI22D1 U1044 ( .A1(n2272), .A2(n973), .B1(n2280), .B2(n2271), .ZN(
        dp_cluster_1_mult_512_C418_n353) );
  OAI22D1 U1045 ( .A1(n2256), .A2(n972), .B1(n2262), .B2(n2255), .ZN(
        dp_cluster_1_mult_512_C418_n339) );
  OAI22D1 U1046 ( .A1(n2240), .A2(n974), .B1(n2244), .B2(n2239), .ZN(
        dp_cluster_1_mult_512_C418_n325) );
  FA1D0 U1047 ( .A(dp_cluster_3_mult_512_C415_n325), .B(
        dp_cluster_3_mult_512_C415_n339), .CI(dp_cluster_3_mult_512_C415_n353), 
        .CO(dp_cluster_3_mult_512_C415_n218), .S(
        dp_cluster_3_mult_512_C415_n219) );
  OAI22D1 U1048 ( .A1(n2923), .A2(n997), .B1(n2931), .B2(n2922), .ZN(
        dp_cluster_3_mult_512_C415_n353) );
  OAI22D1 U1049 ( .A1(n2907), .A2(n996), .B1(n2913), .B2(n2906), .ZN(
        dp_cluster_3_mult_512_C415_n339) );
  OAI22D1 U1050 ( .A1(n2891), .A2(n998), .B1(n2895), .B2(n2890), .ZN(
        dp_cluster_3_mult_512_C415_n325) );
  OAI22D1 U1051 ( .A1(n2216), .A2(n976), .B1(n2304), .B2(n2215), .ZN(
        dp_cluster_1_mult_512_C418_n300) );
  OAI22D1 U1052 ( .A1(n2204), .A2(n971), .B1(n2300), .B2(n2203), .ZN(
        dp_cluster_1_mult_512_C418_n286) );
  OAI22D1 U1053 ( .A1(n2180), .A2(n2306), .B1(n2307), .B2(n2179), .ZN(
        dp_cluster_1_mult_512_C418_n259) );
  OAI22D1 U1054 ( .A1(n2064), .A2(n970), .B1(n2152), .B2(n2063), .ZN(
        dp_cluster_1_mult_513_C418_n300) );
  OAI22D1 U1055 ( .A1(n2052), .A2(n965), .B1(n2148), .B2(n2051), .ZN(
        dp_cluster_1_mult_513_C418_n286) );
  OAI22D1 U1056 ( .A1(n2028), .A2(n2154), .B1(n2155), .B2(n2027), .ZN(
        dp_cluster_1_mult_513_C418_n259) );
  OAI22D1 U1057 ( .A1(n2867), .A2(n1000), .B1(n2955), .B2(n2866), .ZN(
        dp_cluster_3_mult_512_C415_n300) );
  OAI22D1 U1058 ( .A1(n2855), .A2(n995), .B1(n2951), .B2(n2854), .ZN(
        dp_cluster_3_mult_512_C415_n286) );
  OAI22D1 U1059 ( .A1(n2831), .A2(n2957), .B1(n2958), .B2(n2830), .ZN(
        dp_cluster_3_mult_512_C415_n259) );
  OAI22D1 U1060 ( .A1(n2715), .A2(n994), .B1(n2803), .B2(n2714), .ZN(
        dp_cluster_3_mult_513_C415_n300) );
  OAI22D1 U1061 ( .A1(n2703), .A2(n989), .B1(n2799), .B2(n2702), .ZN(
        dp_cluster_3_mult_513_C415_n286) );
  OAI22D1 U1062 ( .A1(n2679), .A2(n2805), .B1(n2806), .B2(n2678), .ZN(
        dp_cluster_3_mult_513_C415_n259) );
  FA1D0 U1063 ( .A(dp_cluster_1_mult_512_C418_n307), .B(
        dp_cluster_1_mult_512_C418_n280), .CI(dp_cluster_1_mult_512_C418_n293), 
        .CO(dp_cluster_1_mult_512_C418_n199), .S(
        dp_cluster_1_mult_512_C418_n200) );
  OAI22D1 U1064 ( .A1(n2223), .A2(n976), .B1(n2304), .B2(n2222), .ZN(
        dp_cluster_1_mult_512_C418_n307) );
  NR2D1 U1065 ( .A1(n2310), .A2(n1098), .ZN(dp_cluster_1_mult_512_C418_n280)
         );
  OAI22D1 U1066 ( .A1(n2211), .A2(n971), .B1(n2300), .B2(n2210), .ZN(
        dp_cluster_1_mult_512_C418_n293) );
  FA1D0 U1067 ( .A(dp_cluster_1_mult_513_C418_n307), .B(
        dp_cluster_1_mult_513_C418_n280), .CI(dp_cluster_1_mult_513_C418_n293), 
        .CO(dp_cluster_1_mult_513_C418_n199), .S(
        dp_cluster_1_mult_513_C418_n200) );
  OAI22D1 U1068 ( .A1(n2071), .A2(n970), .B1(n2152), .B2(n2070), .ZN(
        dp_cluster_1_mult_513_C418_n307) );
  NR2D1 U1069 ( .A1(n2158), .A2(n1092), .ZN(dp_cluster_1_mult_513_C418_n280)
         );
  OAI22D1 U1070 ( .A1(n2059), .A2(n965), .B1(n2148), .B2(n2058), .ZN(
        dp_cluster_1_mult_513_C418_n293) );
  FA1D0 U1071 ( .A(dp_cluster_0_mult_486_C412_n307), .B(
        dp_cluster_0_mult_486_C412_n280), .CI(dp_cluster_0_mult_486_C412_n293), 
        .CO(dp_cluster_0_mult_486_C412_n199), .S(
        dp_cluster_0_mult_486_C412_n200) );
  OAI22D1 U1072 ( .A1(n1745), .A2(n958), .B1(n1826), .B2(n1744), .ZN(
        dp_cluster_0_mult_486_C412_n307) );
  NR2D1 U1073 ( .A1(n1832), .A2(n1100), .ZN(dp_cluster_0_mult_486_C412_n280)
         );
  OAI22D1 U1074 ( .A1(n1733), .A2(n953), .B1(n1822), .B2(n1732), .ZN(
        dp_cluster_0_mult_486_C412_n293) );
  FA1D0 U1075 ( .A(dp_cluster_0_mult_485_C412_n307), .B(
        dp_cluster_0_mult_485_C412_n280), .CI(dp_cluster_0_mult_485_C412_n293), 
        .CO(dp_cluster_0_mult_485_C412_n199), .S(
        dp_cluster_0_mult_485_C412_n200) );
  OAI22D1 U1076 ( .A1(n1897), .A2(n964), .B1(n1978), .B2(n1896), .ZN(
        dp_cluster_0_mult_485_C412_n307) );
  NR2D1 U1077 ( .A1(n1984), .A2(n1094), .ZN(dp_cluster_0_mult_485_C412_n280)
         );
  OAI22D1 U1078 ( .A1(n1885), .A2(n959), .B1(n1974), .B2(n1884), .ZN(
        dp_cluster_0_mult_485_C412_n293) );
  FA1D0 U1079 ( .A(dp_cluster_3_mult_512_C415_n307), .B(
        dp_cluster_3_mult_512_C415_n280), .CI(dp_cluster_3_mult_512_C415_n293), 
        .CO(dp_cluster_3_mult_512_C415_n199), .S(
        dp_cluster_3_mult_512_C415_n200) );
  OAI22D1 U1080 ( .A1(n2874), .A2(n1000), .B1(n2955), .B2(n2873), .ZN(
        dp_cluster_3_mult_512_C415_n307) );
  NR2D1 U1081 ( .A1(n2961), .A2(n1095), .ZN(dp_cluster_3_mult_512_C415_n280)
         );
  OAI22D1 U1082 ( .A1(n2862), .A2(n995), .B1(n2951), .B2(n2861), .ZN(
        dp_cluster_3_mult_512_C415_n293) );
  FA1D0 U1083 ( .A(dp_cluster_3_mult_513_C415_n307), .B(
        dp_cluster_3_mult_513_C415_n280), .CI(dp_cluster_3_mult_513_C415_n293), 
        .CO(dp_cluster_3_mult_513_C415_n199), .S(
        dp_cluster_3_mult_513_C415_n200) );
  OAI22D1 U1084 ( .A1(n2722), .A2(n994), .B1(n2803), .B2(n2721), .ZN(
        dp_cluster_3_mult_513_C415_n307) );
  NR2D1 U1085 ( .A1(n2809), .A2(n1089), .ZN(dp_cluster_3_mult_513_C415_n280)
         );
  OAI22D1 U1086 ( .A1(n2710), .A2(n989), .B1(n2799), .B2(n2709), .ZN(
        dp_cluster_3_mult_513_C415_n293) );
  FA1D0 U1087 ( .A(dp_cluster_2_mult_486_C409_n307), .B(
        dp_cluster_2_mult_486_C409_n280), .CI(dp_cluster_2_mult_486_C409_n293), 
        .CO(dp_cluster_2_mult_486_C409_n199), .S(
        dp_cluster_2_mult_486_C409_n200) );
  OAI22D1 U1088 ( .A1(n2396), .A2(n982), .B1(n2477), .B2(n2395), .ZN(
        dp_cluster_2_mult_486_C409_n307) );
  NR2D1 U1089 ( .A1(n2483), .A2(n1097), .ZN(dp_cluster_2_mult_486_C409_n280)
         );
  OAI22D1 U1090 ( .A1(n2384), .A2(n977), .B1(n2473), .B2(n2383), .ZN(
        dp_cluster_2_mult_486_C409_n293) );
  FA1D0 U1091 ( .A(dp_cluster_2_mult_485_C409_n307), .B(
        dp_cluster_2_mult_485_C409_n280), .CI(dp_cluster_2_mult_485_C409_n293), 
        .CO(dp_cluster_2_mult_485_C409_n199), .S(
        dp_cluster_2_mult_485_C409_n200) );
  OAI22D1 U1092 ( .A1(n2548), .A2(n988), .B1(n2629), .B2(n2547), .ZN(
        dp_cluster_2_mult_485_C409_n307) );
  NR2D1 U1093 ( .A1(n2635), .A2(n1091), .ZN(dp_cluster_2_mult_485_C409_n280)
         );
  OAI22D1 U1094 ( .A1(n2536), .A2(n983), .B1(n2625), .B2(n2535), .ZN(
        dp_cluster_2_mult_485_C409_n293) );
  OAI22D1 U1095 ( .A1(n2224), .A2(n976), .B1(n2304), .B2(n2223), .ZN(
        dp_cluster_1_mult_512_C418_n308) );
  OAI22D1 U1096 ( .A1(n2072), .A2(n970), .B1(n2152), .B2(n2071), .ZN(
        dp_cluster_1_mult_513_C418_n308) );
  OAI22D1 U1097 ( .A1(n1898), .A2(n964), .B1(n1978), .B2(n1897), .ZN(
        dp_cluster_0_mult_485_C412_n308) );
  OAI22D1 U1098 ( .A1(n2875), .A2(n1000), .B1(n2955), .B2(n2874), .ZN(
        dp_cluster_3_mult_512_C415_n308) );
  OAI22D1 U1099 ( .A1(n2723), .A2(n994), .B1(n2803), .B2(n2722), .ZN(
        dp_cluster_3_mult_513_C415_n308) );
  OAI22D1 U1100 ( .A1(n2549), .A2(n988), .B1(n2629), .B2(n2548), .ZN(
        dp_cluster_2_mult_485_C409_n308) );
  OAI22D1 U1101 ( .A1(n1746), .A2(n958), .B1(n1826), .B2(n1745), .ZN(
        dp_cluster_0_mult_486_C412_n308) );
  OAI22D1 U1102 ( .A1(n2397), .A2(n982), .B1(n2477), .B2(n2396), .ZN(
        dp_cluster_2_mult_486_C409_n308) );
  OAI22D1 U1103 ( .A1(n2205), .A2(n971), .B1(n2300), .B2(n2204), .ZN(
        dp_cluster_1_mult_512_C418_n287) );
  OAI22D1 U1104 ( .A1(n2053), .A2(n965), .B1(n2148), .B2(n2052), .ZN(
        dp_cluster_1_mult_513_C418_n287) );
  OAI22D1 U1105 ( .A1(n1727), .A2(n953), .B1(n1822), .B2(n1726), .ZN(
        dp_cluster_0_mult_486_C412_n287) );
  OAI22D1 U1106 ( .A1(n1879), .A2(n959), .B1(n1974), .B2(n1878), .ZN(
        dp_cluster_0_mult_485_C412_n287) );
  OAI22D1 U1107 ( .A1(n2856), .A2(n995), .B1(n2951), .B2(n2855), .ZN(
        dp_cluster_3_mult_512_C415_n287) );
  OAI22D1 U1108 ( .A1(n2704), .A2(n989), .B1(n2799), .B2(n2703), .ZN(
        dp_cluster_3_mult_513_C415_n287) );
  OAI22D1 U1109 ( .A1(n2378), .A2(n977), .B1(n2473), .B2(n2377), .ZN(
        dp_cluster_2_mult_486_C409_n287) );
  OAI22D1 U1110 ( .A1(n2530), .A2(n983), .B1(n2625), .B2(n2529), .ZN(
        dp_cluster_2_mult_485_C409_n287) );
  OAI22D1 U1111 ( .A1(n1757), .A2(n956), .B1(n1766), .B2(n1756), .ZN(
        dp_cluster_0_mult_486_C412_n320) );
  OAI22D1 U1112 ( .A1(n1909), .A2(n962), .B1(n1918), .B2(n1908), .ZN(
        dp_cluster_0_mult_485_C412_n320) );
  OAI22D1 U1113 ( .A1(n2408), .A2(n980), .B1(n2417), .B2(n2407), .ZN(
        dp_cluster_2_mult_486_C409_n320) );
  OAI22D1 U1114 ( .A1(n2560), .A2(n986), .B1(n2569), .B2(n2559), .ZN(
        dp_cluster_2_mult_485_C409_n320) );
  OAI22D1 U1115 ( .A1(n2235), .A2(n974), .B1(n2244), .B2(n2234), .ZN(
        dp_cluster_1_mult_512_C418_n320) );
  OAI22D1 U1116 ( .A1(n2083), .A2(n968), .B1(n2092), .B2(n2082), .ZN(
        dp_cluster_1_mult_513_C418_n320) );
  OAI22D1 U1117 ( .A1(n2886), .A2(n998), .B1(n2895), .B2(n2885), .ZN(
        dp_cluster_3_mult_512_C415_n320) );
  OAI22D1 U1118 ( .A1(n2734), .A2(n992), .B1(n2743), .B2(n2733), .ZN(
        dp_cluster_3_mult_513_C415_n320) );
  OAI22D1 U1119 ( .A1(n2191), .A2(n975), .B1(n2310), .B2(n2190), .ZN(
        dp_cluster_1_mult_512_C418_n272) );
  OAI22D1 U1120 ( .A1(n2039), .A2(n969), .B1(n2158), .B2(n2038), .ZN(
        dp_cluster_1_mult_513_C418_n272) );
  OAI22D1 U1121 ( .A1(n1713), .A2(n957), .B1(n1832), .B2(n1712), .ZN(
        dp_cluster_0_mult_486_C412_n272) );
  OAI22D1 U1122 ( .A1(n1865), .A2(n963), .B1(n1984), .B2(n1864), .ZN(
        dp_cluster_0_mult_485_C412_n272) );
  OAI22D1 U1123 ( .A1(n2842), .A2(n999), .B1(n2961), .B2(n2841), .ZN(
        dp_cluster_3_mult_512_C415_n272) );
  OAI22D1 U1124 ( .A1(n2690), .A2(n993), .B1(n2809), .B2(n2689), .ZN(
        dp_cluster_3_mult_513_C415_n272) );
  OAI22D1 U1125 ( .A1(n2364), .A2(n981), .B1(n2483), .B2(n2363), .ZN(
        dp_cluster_2_mult_486_C409_n272) );
  OAI22D1 U1126 ( .A1(n2516), .A2(n987), .B1(n2635), .B2(n2515), .ZN(
        dp_cluster_2_mult_485_C409_n272) );
  OAI22D1 U1127 ( .A1(n1704), .A2(n1828), .B1(n1829), .B2(n1703), .ZN(
        dp_cluster_0_mult_486_C412_n261) );
  OAI22D1 U1128 ( .A1(n1856), .A2(n1980), .B1(n1981), .B2(n1855), .ZN(
        dp_cluster_0_mult_485_C412_n261) );
  OAI22D1 U1129 ( .A1(n2355), .A2(n2479), .B1(n2480), .B2(n2354), .ZN(
        dp_cluster_2_mult_486_C409_n261) );
  OAI22D1 U1130 ( .A1(n2507), .A2(n2631), .B1(n2632), .B2(n2506), .ZN(
        dp_cluster_2_mult_485_C409_n261) );
  OAI22D1 U1131 ( .A1(n2182), .A2(n2306), .B1(n2307), .B2(n2181), .ZN(
        dp_cluster_1_mult_512_C418_n261) );
  OAI22D1 U1132 ( .A1(n2030), .A2(n2154), .B1(n2155), .B2(n2029), .ZN(
        dp_cluster_1_mult_513_C418_n261) );
  OAI22D1 U1133 ( .A1(n2833), .A2(n2957), .B1(n2958), .B2(n2832), .ZN(
        dp_cluster_3_mult_512_C415_n261) );
  OAI22D1 U1134 ( .A1(n2681), .A2(n2805), .B1(n2806), .B2(n2680), .ZN(
        dp_cluster_3_mult_513_C415_n261) );
  OAI22D1 U1135 ( .A1(n2220), .A2(n976), .B1(n2304), .B2(n2219), .ZN(
        dp_cluster_1_mult_512_C418_n304) );
  OAI22D1 U1136 ( .A1(n2068), .A2(n970), .B1(n2152), .B2(n2067), .ZN(
        dp_cluster_1_mult_513_C418_n304) );
  OAI22D1 U1137 ( .A1(n1742), .A2(n958), .B1(n1826), .B2(n1741), .ZN(
        dp_cluster_0_mult_486_C412_n304) );
  OAI22D1 U1138 ( .A1(n1894), .A2(n964), .B1(n1978), .B2(n1893), .ZN(
        dp_cluster_0_mult_485_C412_n304) );
  OAI22D1 U1139 ( .A1(n2871), .A2(n1000), .B1(n2955), .B2(n2870), .ZN(
        dp_cluster_3_mult_512_C415_n304) );
  OAI22D1 U1140 ( .A1(n2719), .A2(n994), .B1(n2803), .B2(n2718), .ZN(
        dp_cluster_3_mult_513_C415_n304) );
  OAI22D1 U1141 ( .A1(n2393), .A2(n982), .B1(n2477), .B2(n2392), .ZN(
        dp_cluster_2_mult_486_C409_n304) );
  OAI22D1 U1142 ( .A1(n2545), .A2(n988), .B1(n2629), .B2(n2544), .ZN(
        dp_cluster_2_mult_485_C409_n304) );
  OAI22D1 U1143 ( .A1(n2194), .A2(n975), .B1(n2310), .B2(n2193), .ZN(
        dp_cluster_1_mult_512_C418_n275) );
  OAI22D1 U1144 ( .A1(n2042), .A2(n969), .B1(n2158), .B2(n2041), .ZN(
        dp_cluster_1_mult_513_C418_n275) );
  OAI22D1 U1145 ( .A1(n1716), .A2(n957), .B1(n1832), .B2(n1715), .ZN(
        dp_cluster_0_mult_486_C412_n275) );
  OAI22D1 U1146 ( .A1(n1868), .A2(n963), .B1(n1984), .B2(n1867), .ZN(
        dp_cluster_0_mult_485_C412_n275) );
  OAI22D1 U1147 ( .A1(n2845), .A2(n999), .B1(n2961), .B2(n2844), .ZN(
        dp_cluster_3_mult_512_C415_n275) );
  OAI22D1 U1148 ( .A1(n2693), .A2(n993), .B1(n2809), .B2(n2692), .ZN(
        dp_cluster_3_mult_513_C415_n275) );
  OAI22D1 U1149 ( .A1(n2367), .A2(n981), .B1(n2483), .B2(n2366), .ZN(
        dp_cluster_2_mult_486_C409_n275) );
  OAI22D1 U1150 ( .A1(n2519), .A2(n987), .B1(n2635), .B2(n2518), .ZN(
        dp_cluster_2_mult_485_C409_n275) );
  OAI22D1 U1151 ( .A1(n2190), .A2(n975), .B1(n2310), .B2(n2189), .ZN(
        dp_cluster_1_mult_512_C418_n271) );
  OAI22D1 U1152 ( .A1(n2038), .A2(n969), .B1(n2158), .B2(n2037), .ZN(
        dp_cluster_1_mult_513_C418_n271) );
  OAI22D1 U1153 ( .A1(n1712), .A2(n957), .B1(n1832), .B2(n1711), .ZN(
        dp_cluster_0_mult_486_C412_n271) );
  OAI22D1 U1154 ( .A1(n1864), .A2(n963), .B1(n1984), .B2(n1863), .ZN(
        dp_cluster_0_mult_485_C412_n271) );
  OAI22D1 U1155 ( .A1(n2841), .A2(n999), .B1(n2961), .B2(n2840), .ZN(
        dp_cluster_3_mult_512_C415_n271) );
  OAI22D1 U1156 ( .A1(n2689), .A2(n993), .B1(n2809), .B2(n2688), .ZN(
        dp_cluster_3_mult_513_C415_n271) );
  OAI22D1 U1157 ( .A1(n2363), .A2(n981), .B1(n2483), .B2(n2362), .ZN(
        dp_cluster_2_mult_486_C409_n271) );
  OAI22D1 U1158 ( .A1(n2515), .A2(n987), .B1(n2635), .B2(n2514), .ZN(
        dp_cluster_2_mult_485_C409_n271) );
  OAI22D1 U1159 ( .A1(n1699), .A2(n1828), .B1(n1829), .B2(n1698), .ZN(
        dp_cluster_0_mult_486_C412_n256) );
  OAI22D1 U1160 ( .A1(n1851), .A2(n1980), .B1(n1981), .B2(n1850), .ZN(
        dp_cluster_0_mult_485_C412_n256) );
  OAI22D1 U1161 ( .A1(n2350), .A2(n2479), .B1(n2480), .B2(n2349), .ZN(
        dp_cluster_2_mult_486_C409_n256) );
  OAI22D1 U1162 ( .A1(n2502), .A2(n2631), .B1(n2632), .B2(n2501), .ZN(
        dp_cluster_2_mult_485_C409_n256) );
  OAI22D1 U1163 ( .A1(n2177), .A2(n2306), .B1(n2307), .B2(n2176), .ZN(
        dp_cluster_1_mult_512_C418_n256) );
  OAI22D1 U1164 ( .A1(n2025), .A2(n2154), .B1(n2155), .B2(n2024), .ZN(
        dp_cluster_1_mult_513_C418_n256) );
  OAI22D1 U1165 ( .A1(n2828), .A2(n2957), .B1(n2958), .B2(n2827), .ZN(
        dp_cluster_3_mult_512_C415_n256) );
  OAI22D1 U1166 ( .A1(n2676), .A2(n2805), .B1(n2806), .B2(n2675), .ZN(
        dp_cluster_3_mult_513_C415_n256) );
  OAI22D1 U1167 ( .A1(n1933), .A2(n960), .B1(n1936), .B2(n1932), .ZN(
        dp_cluster_0_mult_485_C412_n342) );
  OAI22D1 U1168 ( .A1(n2584), .A2(n984), .B1(n2587), .B2(n2583), .ZN(
        dp_cluster_2_mult_485_C409_n342) );
  OAI22D1 U1169 ( .A1(n2225), .A2(n976), .B1(n2304), .B2(n2224), .ZN(
        dp_cluster_1_mult_512_C418_n309) );
  OAI22D1 U1170 ( .A1(n2073), .A2(n970), .B1(n2152), .B2(n2072), .ZN(
        dp_cluster_1_mult_513_C418_n309) );
  OAI22D1 U1171 ( .A1(n1899), .A2(n964), .B1(n1978), .B2(n1898), .ZN(
        dp_cluster_0_mult_485_C412_n309) );
  OAI22D1 U1172 ( .A1(n2876), .A2(n1000), .B1(n2955), .B2(n2875), .ZN(
        dp_cluster_3_mult_512_C415_n309) );
  OAI22D1 U1173 ( .A1(n2724), .A2(n994), .B1(n2803), .B2(n2723), .ZN(
        dp_cluster_3_mult_513_C415_n309) );
  OAI22D1 U1174 ( .A1(n2550), .A2(n988), .B1(n2629), .B2(n2549), .ZN(
        dp_cluster_2_mult_485_C409_n309) );
  OAI22D1 U1175 ( .A1(n2107), .A2(n966), .B1(n2110), .B2(n2106), .ZN(
        dp_cluster_1_mult_513_C418_n342) );
  OAI22D1 U1176 ( .A1(n2758), .A2(n990), .B1(n2761), .B2(n2757), .ZN(
        dp_cluster_3_mult_513_C415_n342) );
  OAI22D1 U1177 ( .A1(n2259), .A2(n972), .B1(n2262), .B2(n2258), .ZN(
        dp_cluster_1_mult_512_C418_n342) );
  OAI22D1 U1178 ( .A1(n2910), .A2(n996), .B1(n2913), .B2(n2909), .ZN(
        dp_cluster_3_mult_512_C415_n342) );
  OAI22D1 U1179 ( .A1(n1781), .A2(n954), .B1(n1784), .B2(n1780), .ZN(
        dp_cluster_0_mult_486_C412_n342) );
  OAI22D1 U1180 ( .A1(n2432), .A2(n978), .B1(n2435), .B2(n2431), .ZN(
        dp_cluster_2_mult_486_C409_n342) );
  OAI22D1 U1181 ( .A1(n1747), .A2(n958), .B1(n1826), .B2(n1746), .ZN(
        dp_cluster_0_mult_486_C412_n309) );
  OAI22D1 U1182 ( .A1(n2398), .A2(n982), .B1(n2477), .B2(n2397), .ZN(
        dp_cluster_2_mult_486_C409_n309) );
  OAI22D1 U1183 ( .A1(n2197), .A2(n975), .B1(n2310), .B2(n2196), .ZN(
        dp_cluster_1_mult_512_C418_n278) );
  OAI22D1 U1184 ( .A1(n2045), .A2(n969), .B1(n2158), .B2(n2044), .ZN(
        dp_cluster_1_mult_513_C418_n278) );
  OAI22D1 U1185 ( .A1(n1719), .A2(n957), .B1(n1832), .B2(n1718), .ZN(
        dp_cluster_0_mult_486_C412_n278) );
  OAI22D1 U1186 ( .A1(n1871), .A2(n963), .B1(n1984), .B2(n1870), .ZN(
        dp_cluster_0_mult_485_C412_n278) );
  OAI22D1 U1187 ( .A1(n2848), .A2(n999), .B1(n2961), .B2(n2847), .ZN(
        dp_cluster_3_mult_512_C415_n278) );
  OAI22D1 U1188 ( .A1(n2696), .A2(n993), .B1(n2809), .B2(n2695), .ZN(
        dp_cluster_3_mult_513_C415_n278) );
  OAI22D1 U1189 ( .A1(n2370), .A2(n981), .B1(n2483), .B2(n2369), .ZN(
        dp_cluster_2_mult_486_C409_n278) );
  OAI22D1 U1190 ( .A1(n2522), .A2(n987), .B1(n2635), .B2(n2521), .ZN(
        dp_cluster_2_mult_485_C409_n278) );
  ND2D1 U1191 ( .A1(n1107), .A2(n1042), .ZN(n1970) );
  ND2D1 U1192 ( .A1(n1110), .A2(n1020), .ZN(n2621) );
  ND2D1 U1193 ( .A1(n1101), .A2(n1086), .ZN(n2144) );
  ND2D1 U1194 ( .A1(n1104), .A2(n1064), .ZN(n2795) );
  ND2D1 U1195 ( .A1(n1107), .A2(n1042), .ZN(n2296) );
  ND2D1 U1196 ( .A1(n1101), .A2(n1086), .ZN(n1818) );
  ND2D1 U1197 ( .A1(n1110), .A2(n1020), .ZN(n2947) );
  ND2D1 U1198 ( .A1(n1104), .A2(n1064), .ZN(n2469) );
  OA22D0 U1199 ( .A1(n2195), .A2(n975), .B1(n2310), .B2(n2194), .Z(n2170) );
  OA22D0 U1200 ( .A1(n2043), .A2(n969), .B1(n2158), .B2(n2042), .Z(n2018) );
  OA22D0 U1201 ( .A1(n1717), .A2(n957), .B1(n1832), .B2(n1716), .Z(n1692) );
  OA22D0 U1202 ( .A1(n1869), .A2(n963), .B1(n1984), .B2(n1868), .Z(n1844) );
  OA22D0 U1203 ( .A1(n2846), .A2(n999), .B1(n2961), .B2(n2845), .Z(n2821) );
  OA22D0 U1204 ( .A1(n2694), .A2(n993), .B1(n2809), .B2(n2693), .Z(n2669) );
  OA22D0 U1205 ( .A1(n2368), .A2(n981), .B1(n2483), .B2(n2367), .Z(n2343) );
  OA22D0 U1206 ( .A1(n2520), .A2(n987), .B1(n2635), .B2(n2519), .Z(n2495) );
  OA22D0 U1207 ( .A1(n2233), .A2(n974), .B1(n2244), .B2(n2232), .Z(n2169) );
  OA22D0 U1208 ( .A1(n2081), .A2(n968), .B1(n2092), .B2(n2080), .Z(n2017) );
  OA22D0 U1209 ( .A1(n2884), .A2(n998), .B1(n2895), .B2(n2883), .Z(n2820) );
  OA22D0 U1210 ( .A1(n2732), .A2(n992), .B1(n2743), .B2(n2731), .Z(n2668) );
  OA22D0 U1211 ( .A1(n1755), .A2(n956), .B1(n1766), .B2(n1754), .Z(n1691) );
  OA22D0 U1212 ( .A1(n1907), .A2(n962), .B1(n1918), .B2(n1906), .Z(n1843) );
  OA22D0 U1213 ( .A1(n2406), .A2(n980), .B1(n2417), .B2(n2405), .Z(n2342) );
  OA22D0 U1214 ( .A1(n2558), .A2(n986), .B1(n2569), .B2(n2557), .Z(n2494) );
  OAI22D1 U1215 ( .A1(n2253), .A2(n972), .B1(n2262), .B2(n2252), .ZN(
        dp_cluster_1_mult_512_C418_n336) );
  OAI22D1 U1216 ( .A1(n2101), .A2(n966), .B1(n2110), .B2(n2100), .ZN(
        dp_cluster_1_mult_513_C418_n336) );
  OAI22D1 U1217 ( .A1(n1775), .A2(n954), .B1(n1784), .B2(n1774), .ZN(
        dp_cluster_0_mult_486_C412_n336) );
  OAI22D1 U1218 ( .A1(n1927), .A2(n960), .B1(n1936), .B2(n1926), .ZN(
        dp_cluster_0_mult_485_C412_n336) );
  OAI22D1 U1219 ( .A1(n2904), .A2(n996), .B1(n2913), .B2(n2903), .ZN(
        dp_cluster_3_mult_512_C415_n336) );
  OAI22D1 U1220 ( .A1(n2752), .A2(n990), .B1(n2761), .B2(n2751), .ZN(
        dp_cluster_3_mult_513_C415_n336) );
  OAI22D1 U1221 ( .A1(n2426), .A2(n978), .B1(n2435), .B2(n2425), .ZN(
        dp_cluster_2_mult_486_C409_n336) );
  OAI22D1 U1222 ( .A1(n2578), .A2(n984), .B1(n2587), .B2(n2577), .ZN(
        dp_cluster_2_mult_485_C409_n336) );
  INVD1 U1223 ( .I(dp_cluster_1_mult_512_C418_n150), .ZN(n1172) );
  OAI22D1 U1224 ( .A1(n2248), .A2(n972), .B1(n2262), .B2(n2247), .ZN(
        dp_cluster_1_mult_512_C418_n331) );
  ND2D1 U1225 ( .A1(n2169), .A2(n2170), .ZN(dp_cluster_1_mult_512_C418_n161)
         );
  INVD1 U1226 ( .I(dp_cluster_1_mult_513_C418_n150), .ZN(n1303) );
  OAI22D1 U1227 ( .A1(n2096), .A2(n966), .B1(n2110), .B2(n2095), .ZN(
        dp_cluster_1_mult_513_C418_n331) );
  ND2D1 U1228 ( .A1(n2017), .A2(n2018), .ZN(dp_cluster_1_mult_513_C418_n161)
         );
  INVD1 U1229 ( .I(dp_cluster_0_mult_486_C412_n150), .ZN(n1302) );
  OAI22D1 U1230 ( .A1(n1770), .A2(n954), .B1(n1784), .B2(n1769), .ZN(
        dp_cluster_0_mult_486_C412_n331) );
  ND2D1 U1231 ( .A1(n1691), .A2(n1692), .ZN(dp_cluster_0_mult_486_C412_n161)
         );
  INVD1 U1232 ( .I(dp_cluster_0_mult_485_C412_n150), .ZN(n1170) );
  OAI22D1 U1233 ( .A1(n1922), .A2(n960), .B1(n1936), .B2(n1921), .ZN(
        dp_cluster_0_mult_485_C412_n331) );
  ND2D1 U1234 ( .A1(n1843), .A2(n1844), .ZN(dp_cluster_0_mult_485_C412_n161)
         );
  INVD1 U1235 ( .I(dp_cluster_3_mult_512_C415_n150), .ZN(n1133) );
  OAI22D1 U1236 ( .A1(n2899), .A2(n996), .B1(n2913), .B2(n2898), .ZN(
        dp_cluster_3_mult_512_C415_n331) );
  ND2D1 U1237 ( .A1(n2820), .A2(n2821), .ZN(dp_cluster_3_mult_512_C415_n161)
         );
  INVD1 U1238 ( .I(dp_cluster_3_mult_513_C415_n150), .ZN(n1270) );
  OAI22D1 U1239 ( .A1(n2747), .A2(n990), .B1(n2761), .B2(n2746), .ZN(
        dp_cluster_3_mult_513_C415_n331) );
  ND2D1 U1240 ( .A1(n2668), .A2(n2669), .ZN(dp_cluster_3_mult_513_C415_n161)
         );
  INVD1 U1241 ( .I(dp_cluster_2_mult_486_C409_n150), .ZN(n1269) );
  OAI22D1 U1242 ( .A1(n2421), .A2(n978), .B1(n2435), .B2(n2420), .ZN(
        dp_cluster_2_mult_486_C409_n331) );
  ND2D1 U1243 ( .A1(n2342), .A2(n2343), .ZN(dp_cluster_2_mult_486_C409_n161)
         );
  INVD1 U1244 ( .I(dp_cluster_2_mult_485_C409_n150), .ZN(n1131) );
  OAI22D1 U1245 ( .A1(n2573), .A2(n984), .B1(n2587), .B2(n2572), .ZN(
        dp_cluster_2_mult_485_C409_n331) );
  ND2D1 U1246 ( .A1(n2494), .A2(n2495), .ZN(dp_cluster_2_mult_485_C409_n161)
         );
  OAI22D1 U1247 ( .A1(n2265), .A2(n973), .B1(n2280), .B2(n2264), .ZN(
        dp_cluster_1_mult_512_C418_n346) );
  OAI22D1 U1248 ( .A1(n2249), .A2(n972), .B1(n2262), .B2(n2248), .ZN(
        dp_cluster_1_mult_512_C418_n332) );
  OAI22D1 U1249 ( .A1(n2219), .A2(n976), .B1(n2304), .B2(n2218), .ZN(
        dp_cluster_1_mult_512_C418_n303) );
  OAI22D1 U1250 ( .A1(n2113), .A2(n967), .B1(n2128), .B2(n2112), .ZN(
        dp_cluster_1_mult_513_C418_n346) );
  OAI22D1 U1251 ( .A1(n2097), .A2(n966), .B1(n2110), .B2(n2096), .ZN(
        dp_cluster_1_mult_513_C418_n332) );
  OAI22D1 U1252 ( .A1(n2067), .A2(n970), .B1(n2152), .B2(n2066), .ZN(
        dp_cluster_1_mult_513_C418_n303) );
  OAI22D1 U1253 ( .A1(n1787), .A2(n955), .B1(n1802), .B2(n1786), .ZN(
        dp_cluster_0_mult_486_C412_n346) );
  OAI22D1 U1254 ( .A1(n1771), .A2(n954), .B1(n1784), .B2(n1770), .ZN(
        dp_cluster_0_mult_486_C412_n332) );
  OAI22D1 U1255 ( .A1(n1741), .A2(n958), .B1(n1826), .B2(n1740), .ZN(
        dp_cluster_0_mult_486_C412_n303) );
  OAI22D1 U1256 ( .A1(n1939), .A2(n961), .B1(n1954), .B2(n1938), .ZN(
        dp_cluster_0_mult_485_C412_n346) );
  OAI22D1 U1257 ( .A1(n1923), .A2(n960), .B1(n1936), .B2(n1922), .ZN(
        dp_cluster_0_mult_485_C412_n332) );
  OAI22D1 U1258 ( .A1(n1893), .A2(n964), .B1(n1978), .B2(n1892), .ZN(
        dp_cluster_0_mult_485_C412_n303) );
  OAI22D1 U1259 ( .A1(n2916), .A2(n997), .B1(n2931), .B2(n2915), .ZN(
        dp_cluster_3_mult_512_C415_n346) );
  OAI22D1 U1260 ( .A1(n2900), .A2(n996), .B1(n2913), .B2(n2899), .ZN(
        dp_cluster_3_mult_512_C415_n332) );
  OAI22D1 U1261 ( .A1(n2870), .A2(n1000), .B1(n2955), .B2(n2869), .ZN(
        dp_cluster_3_mult_512_C415_n303) );
  OAI22D1 U1262 ( .A1(n2764), .A2(n991), .B1(n2779), .B2(n2763), .ZN(
        dp_cluster_3_mult_513_C415_n346) );
  OAI22D1 U1263 ( .A1(n2748), .A2(n990), .B1(n2761), .B2(n2747), .ZN(
        dp_cluster_3_mult_513_C415_n332) );
  OAI22D1 U1264 ( .A1(n2718), .A2(n994), .B1(n2803), .B2(n2717), .ZN(
        dp_cluster_3_mult_513_C415_n303) );
  OAI22D1 U1265 ( .A1(n2438), .A2(n979), .B1(n2453), .B2(n2437), .ZN(
        dp_cluster_2_mult_486_C409_n346) );
  OAI22D1 U1266 ( .A1(n2422), .A2(n978), .B1(n2435), .B2(n2421), .ZN(
        dp_cluster_2_mult_486_C409_n332) );
  OAI22D1 U1267 ( .A1(n2392), .A2(n982), .B1(n2477), .B2(n2391), .ZN(
        dp_cluster_2_mult_486_C409_n303) );
  OAI22D1 U1268 ( .A1(n2590), .A2(n985), .B1(n2605), .B2(n2589), .ZN(
        dp_cluster_2_mult_485_C409_n346) );
  OAI22D1 U1269 ( .A1(n2574), .A2(n984), .B1(n2587), .B2(n2573), .ZN(
        dp_cluster_2_mult_485_C409_n332) );
  OAI22D1 U1270 ( .A1(n2544), .A2(n988), .B1(n2629), .B2(n2543), .ZN(
        dp_cluster_2_mult_485_C409_n303) );
  OAI22D1 U1271 ( .A1(n1738), .A2(n958), .B1(n1826), .B2(n1737), .ZN(
        dp_cluster_0_mult_486_C412_n300) );
  OAI22D1 U1272 ( .A1(n1726), .A2(n953), .B1(n1822), .B2(n1725), .ZN(
        dp_cluster_0_mult_486_C412_n286) );
  OAI22D1 U1273 ( .A1(n1702), .A2(n1828), .B1(n1829), .B2(n1701), .ZN(
        dp_cluster_0_mult_486_C412_n259) );
  OAI22D1 U1274 ( .A1(n1890), .A2(n964), .B1(n1978), .B2(n1889), .ZN(
        dp_cluster_0_mult_485_C412_n300) );
  OAI22D1 U1275 ( .A1(n1878), .A2(n959), .B1(n1974), .B2(n1877), .ZN(
        dp_cluster_0_mult_485_C412_n286) );
  OAI22D1 U1276 ( .A1(n1854), .A2(n1980), .B1(n1981), .B2(n1853), .ZN(
        dp_cluster_0_mult_485_C412_n259) );
  OAI22D1 U1277 ( .A1(n2389), .A2(n982), .B1(n2477), .B2(n2388), .ZN(
        dp_cluster_2_mult_486_C409_n300) );
  OAI22D1 U1278 ( .A1(n2377), .A2(n977), .B1(n2473), .B2(n2376), .ZN(
        dp_cluster_2_mult_486_C409_n286) );
  OAI22D1 U1279 ( .A1(n2353), .A2(n2479), .B1(n2480), .B2(n2352), .ZN(
        dp_cluster_2_mult_486_C409_n259) );
  OAI22D1 U1280 ( .A1(n2541), .A2(n988), .B1(n2629), .B2(n2540), .ZN(
        dp_cluster_2_mult_485_C409_n300) );
  OAI22D1 U1281 ( .A1(n2529), .A2(n983), .B1(n2625), .B2(n2528), .ZN(
        dp_cluster_2_mult_485_C409_n286) );
  OAI22D1 U1282 ( .A1(n2505), .A2(n2631), .B1(n2632), .B2(n2504), .ZN(
        dp_cluster_2_mult_485_C409_n259) );
  OAI22D1 U1283 ( .A1(n2178), .A2(n2306), .B1(n2307), .B2(n2177), .ZN(
        dp_cluster_1_mult_512_C418_n257) );
  OAI22D1 U1284 ( .A1(n2026), .A2(n2154), .B1(n2155), .B2(n2025), .ZN(
        dp_cluster_1_mult_513_C418_n257) );
  OAI22D1 U1285 ( .A1(n1700), .A2(n1828), .B1(n1829), .B2(n1699), .ZN(
        dp_cluster_0_mult_486_C412_n257) );
  OAI22D1 U1286 ( .A1(n1852), .A2(n1980), .B1(n1981), .B2(n1851), .ZN(
        dp_cluster_0_mult_485_C412_n257) );
  OAI22D1 U1287 ( .A1(n2829), .A2(n2957), .B1(n2958), .B2(n2828), .ZN(
        dp_cluster_3_mult_512_C415_n257) );
  OAI22D1 U1288 ( .A1(n2677), .A2(n2805), .B1(n2806), .B2(n2676), .ZN(
        dp_cluster_3_mult_513_C415_n257) );
  OAI22D1 U1289 ( .A1(n2351), .A2(n2479), .B1(n2480), .B2(n2350), .ZN(
        dp_cluster_2_mult_486_C409_n257) );
  OAI22D1 U1290 ( .A1(n2503), .A2(n2631), .B1(n2632), .B2(n2502), .ZN(
        dp_cluster_2_mult_485_C409_n257) );
  OAI22D1 U1291 ( .A1(n2189), .A2(n975), .B1(n2310), .B2(n2188), .ZN(
        dp_cluster_1_mult_512_C418_n270) );
  OAI22D1 U1292 ( .A1(n2037), .A2(n969), .B1(n2158), .B2(n2036), .ZN(
        dp_cluster_1_mult_513_C418_n270) );
  OAI22D1 U1293 ( .A1(n1711), .A2(n957), .B1(n1832), .B2(n1710), .ZN(
        dp_cluster_0_mult_486_C412_n270) );
  OAI22D1 U1294 ( .A1(n1863), .A2(n963), .B1(n1984), .B2(n1862), .ZN(
        dp_cluster_0_mult_485_C412_n270) );
  OAI22D1 U1295 ( .A1(n2840), .A2(n999), .B1(n2961), .B2(n2839), .ZN(
        dp_cluster_3_mult_512_C415_n270) );
  OAI22D1 U1296 ( .A1(n2688), .A2(n993), .B1(n2809), .B2(n2687), .ZN(
        dp_cluster_3_mult_513_C415_n270) );
  OAI22D1 U1297 ( .A1(n2362), .A2(n981), .B1(n2483), .B2(n2361), .ZN(
        dp_cluster_2_mult_486_C409_n270) );
  OAI22D1 U1298 ( .A1(n2514), .A2(n987), .B1(n2635), .B2(n2513), .ZN(
        dp_cluster_2_mult_485_C409_n270) );
  OAI22D1 U1299 ( .A1(n2200), .A2(n971), .B1(n2300), .B2(n2199), .ZN(
        dp_cluster_1_mult_512_C418_n283) );
  OAI22D1 U1300 ( .A1(n2048), .A2(n965), .B1(n2148), .B2(n2047), .ZN(
        dp_cluster_1_mult_513_C418_n283) );
  OAI22D1 U1301 ( .A1(n1722), .A2(n953), .B1(n1822), .B2(n1721), .ZN(
        dp_cluster_0_mult_486_C412_n283) );
  OAI22D1 U1302 ( .A1(n1874), .A2(n959), .B1(n1974), .B2(n1873), .ZN(
        dp_cluster_0_mult_485_C412_n283) );
  OAI22D1 U1303 ( .A1(n2851), .A2(n995), .B1(n2951), .B2(n2850), .ZN(
        dp_cluster_3_mult_512_C415_n283) );
  OAI22D1 U1304 ( .A1(n2699), .A2(n989), .B1(n2799), .B2(n2698), .ZN(
        dp_cluster_3_mult_513_C415_n283) );
  OAI22D1 U1305 ( .A1(n2373), .A2(n977), .B1(n2473), .B2(n2372), .ZN(
        dp_cluster_2_mult_486_C409_n283) );
  OAI22D1 U1306 ( .A1(n2525), .A2(n983), .B1(n2625), .B2(n2524), .ZN(
        dp_cluster_2_mult_485_C409_n283) );
  INR2D1 U1307 ( .A1(dp_cluster_0_N85), .B1(dp_cluster_0_N57), .ZN(n1991) );
  NR2D1 U1308 ( .A1(n1044), .A2(n1093), .ZN(dp_cluster_0_N57) );
  NR2D1 U1309 ( .A1(n1088), .A2(n1099), .ZN(dp_cluster_0_N85) );
  INR2D1 U1310 ( .A1(dp_cluster_2_N29), .B1(dp_cluster_2_N1), .ZN(n2642) );
  NR2D1 U1311 ( .A1(n1022), .A2(n1090), .ZN(dp_cluster_2_N1) );
  NR2D1 U1312 ( .A1(n1066), .A2(n1096), .ZN(dp_cluster_2_N29) );
  FA1D0 U1313 ( .A(dp_cluster_0_mult_485_C412_n234), .B(
        dp_cluster_0_mult_485_C412_n235), .CI(dp_cluster_0_mult_485_C412_n73), 
        .CO(dp_cluster_0_mult_485_C412_n72), .S(dp_cluster_0_N63) );
  FA1D0 U1314 ( .A(dp_cluster_2_mult_485_C409_n234), .B(
        dp_cluster_2_mult_485_C409_n235), .CI(dp_cluster_2_mult_485_C409_n73), 
        .CO(dp_cluster_2_mult_485_C409_n72), .S(dp_cluster_2_N7) );
  OAI22D1 U1315 ( .A1(n2232), .A2(n974), .B1(n2244), .B2(n2231), .ZN(
        dp_cluster_1_mult_512_C418_n317) );
  OAI22D1 U1316 ( .A1(n2218), .A2(n976), .B1(n2304), .B2(n2217), .ZN(
        dp_cluster_1_mult_512_C418_n302) );
  OAI22D1 U1317 ( .A1(n2206), .A2(n971), .B1(n2300), .B2(n2205), .ZN(
        dp_cluster_1_mult_512_C418_n288) );
  OAI22D1 U1318 ( .A1(n2080), .A2(n968), .B1(n2092), .B2(n2079), .ZN(
        dp_cluster_1_mult_513_C418_n317) );
  OAI22D1 U1319 ( .A1(n2066), .A2(n970), .B1(n2152), .B2(n2065), .ZN(
        dp_cluster_1_mult_513_C418_n302) );
  OAI22D1 U1320 ( .A1(n2054), .A2(n965), .B1(n2148), .B2(n2053), .ZN(
        dp_cluster_1_mult_513_C418_n288) );
  OAI22D1 U1321 ( .A1(n1754), .A2(n956), .B1(n1766), .B2(n1753), .ZN(
        dp_cluster_0_mult_486_C412_n317) );
  OAI22D1 U1322 ( .A1(n1740), .A2(n958), .B1(n1826), .B2(n1739), .ZN(
        dp_cluster_0_mult_486_C412_n302) );
  OAI22D1 U1323 ( .A1(n1728), .A2(n953), .B1(n1822), .B2(n1727), .ZN(
        dp_cluster_0_mult_486_C412_n288) );
  OAI22D1 U1324 ( .A1(n1906), .A2(n962), .B1(n1918), .B2(n1905), .ZN(
        dp_cluster_0_mult_485_C412_n317) );
  OAI22D1 U1325 ( .A1(n1892), .A2(n964), .B1(n1978), .B2(n1891), .ZN(
        dp_cluster_0_mult_485_C412_n302) );
  OAI22D1 U1326 ( .A1(n1880), .A2(n959), .B1(n1974), .B2(n1879), .ZN(
        dp_cluster_0_mult_485_C412_n288) );
  OAI22D1 U1327 ( .A1(n2883), .A2(n998), .B1(n2895), .B2(n2882), .ZN(
        dp_cluster_3_mult_512_C415_n317) );
  OAI22D1 U1328 ( .A1(n2869), .A2(n1000), .B1(n2955), .B2(n2868), .ZN(
        dp_cluster_3_mult_512_C415_n302) );
  OAI22D1 U1329 ( .A1(n2857), .A2(n995), .B1(n2951), .B2(n2856), .ZN(
        dp_cluster_3_mult_512_C415_n288) );
  OAI22D1 U1330 ( .A1(n2731), .A2(n992), .B1(n2743), .B2(n2730), .ZN(
        dp_cluster_3_mult_513_C415_n317) );
  OAI22D1 U1331 ( .A1(n2717), .A2(n994), .B1(n2803), .B2(n2716), .ZN(
        dp_cluster_3_mult_513_C415_n302) );
  OAI22D1 U1332 ( .A1(n2705), .A2(n989), .B1(n2799), .B2(n2704), .ZN(
        dp_cluster_3_mult_513_C415_n288) );
  OAI22D1 U1333 ( .A1(n2405), .A2(n980), .B1(n2417), .B2(n2404), .ZN(
        dp_cluster_2_mult_486_C409_n317) );
  OAI22D1 U1334 ( .A1(n2391), .A2(n982), .B1(n2477), .B2(n2390), .ZN(
        dp_cluster_2_mult_486_C409_n302) );
  OAI22D1 U1335 ( .A1(n2379), .A2(n977), .B1(n2473), .B2(n2378), .ZN(
        dp_cluster_2_mult_486_C409_n288) );
  OAI22D1 U1336 ( .A1(n2557), .A2(n986), .B1(n2569), .B2(n2556), .ZN(
        dp_cluster_2_mult_485_C409_n317) );
  OAI22D1 U1337 ( .A1(n2543), .A2(n988), .B1(n2629), .B2(n2542), .ZN(
        dp_cluster_2_mult_485_C409_n302) );
  OAI22D1 U1338 ( .A1(n2531), .A2(n983), .B1(n2625), .B2(n2530), .ZN(
        dp_cluster_2_mult_485_C409_n288) );
  OAI22D1 U1339 ( .A1(n2247), .A2(n972), .B1(n2262), .B2(n2246), .ZN(
        dp_cluster_1_mult_512_C418_n330) );
  OAI22D1 U1340 ( .A1(n2231), .A2(n974), .B1(n2244), .B2(n2230), .ZN(
        dp_cluster_1_mult_512_C418_n316) );
  OAI22D1 U1341 ( .A1(n2217), .A2(n976), .B1(n2304), .B2(n2216), .ZN(
        dp_cluster_1_mult_512_C418_n301) );
  OAI22D1 U1342 ( .A1(n2095), .A2(n966), .B1(n2110), .B2(n2094), .ZN(
        dp_cluster_1_mult_513_C418_n330) );
  OAI22D1 U1343 ( .A1(n2079), .A2(n968), .B1(n2092), .B2(n2078), .ZN(
        dp_cluster_1_mult_513_C418_n316) );
  OAI22D1 U1344 ( .A1(n2065), .A2(n970), .B1(n2152), .B2(n2064), .ZN(
        dp_cluster_1_mult_513_C418_n301) );
  OAI22D1 U1345 ( .A1(n1769), .A2(n954), .B1(n1784), .B2(n1768), .ZN(
        dp_cluster_0_mult_486_C412_n330) );
  OAI22D1 U1346 ( .A1(n1753), .A2(n956), .B1(n1766), .B2(n1752), .ZN(
        dp_cluster_0_mult_486_C412_n316) );
  OAI22D1 U1347 ( .A1(n1739), .A2(n958), .B1(n1826), .B2(n1738), .ZN(
        dp_cluster_0_mult_486_C412_n301) );
  OAI22D1 U1348 ( .A1(n1921), .A2(n960), .B1(n1936), .B2(n1920), .ZN(
        dp_cluster_0_mult_485_C412_n330) );
  OAI22D1 U1349 ( .A1(n1905), .A2(n962), .B1(n1918), .B2(n1904), .ZN(
        dp_cluster_0_mult_485_C412_n316) );
  OAI22D1 U1350 ( .A1(n1891), .A2(n964), .B1(n1978), .B2(n1890), .ZN(
        dp_cluster_0_mult_485_C412_n301) );
  OAI22D1 U1351 ( .A1(n2898), .A2(n996), .B1(n2913), .B2(n2897), .ZN(
        dp_cluster_3_mult_512_C415_n330) );
  OAI22D1 U1352 ( .A1(n2882), .A2(n998), .B1(n2895), .B2(n2881), .ZN(
        dp_cluster_3_mult_512_C415_n316) );
  OAI22D1 U1353 ( .A1(n2868), .A2(n1000), .B1(n2955), .B2(n2867), .ZN(
        dp_cluster_3_mult_512_C415_n301) );
  OAI22D1 U1354 ( .A1(n2746), .A2(n990), .B1(n2761), .B2(n2745), .ZN(
        dp_cluster_3_mult_513_C415_n330) );
  OAI22D1 U1355 ( .A1(n2730), .A2(n992), .B1(n2743), .B2(n2729), .ZN(
        dp_cluster_3_mult_513_C415_n316) );
  OAI22D1 U1356 ( .A1(n2716), .A2(n994), .B1(n2803), .B2(n2715), .ZN(
        dp_cluster_3_mult_513_C415_n301) );
  OAI22D1 U1357 ( .A1(n2420), .A2(n978), .B1(n2435), .B2(n2419), .ZN(
        dp_cluster_2_mult_486_C409_n330) );
  OAI22D1 U1358 ( .A1(n2404), .A2(n980), .B1(n2417), .B2(n2403), .ZN(
        dp_cluster_2_mult_486_C409_n316) );
  OAI22D1 U1359 ( .A1(n2390), .A2(n982), .B1(n2477), .B2(n2389), .ZN(
        dp_cluster_2_mult_486_C409_n301) );
  OAI22D1 U1360 ( .A1(n2572), .A2(n984), .B1(n2587), .B2(n2571), .ZN(
        dp_cluster_2_mult_485_C409_n330) );
  OAI22D1 U1361 ( .A1(n2556), .A2(n986), .B1(n2569), .B2(n2555), .ZN(
        dp_cluster_2_mult_485_C409_n316) );
  OAI22D1 U1362 ( .A1(n2542), .A2(n988), .B1(n2629), .B2(n2541), .ZN(
        dp_cluster_2_mult_485_C409_n301) );
  XOR3D1 U1363 ( .A1(dp_cluster_1_mult_512_C418_n81), .A2(
        dp_cluster_1_mult_512_C418_n80), .A3(dp_cluster_1_mult_512_C418_n52), 
        .Z(n2314) );
  XOR3D1 U1364 ( .A1(dp_cluster_1_mult_513_C418_n81), .A2(
        dp_cluster_1_mult_513_C418_n80), .A3(dp_cluster_1_mult_513_C418_n52), 
        .Z(n2162) );
  XOR3D1 U1365 ( .A1(dp_cluster_0_mult_485_C412_n81), .A2(
        dp_cluster_0_mult_485_C412_n80), .A3(dp_cluster_0_mult_485_C412_n52), 
        .Z(n1988) );
  XOR3D1 U1366 ( .A1(dp_cluster_3_mult_512_C415_n81), .A2(
        dp_cluster_3_mult_512_C415_n80), .A3(dp_cluster_3_mult_512_C415_n52), 
        .Z(n2965) );
  XOR3D1 U1367 ( .A1(dp_cluster_3_mult_513_C415_n81), .A2(
        dp_cluster_3_mult_513_C415_n80), .A3(dp_cluster_3_mult_513_C415_n52), 
        .Z(n2813) );
  XOR3D1 U1368 ( .A1(dp_cluster_2_mult_485_C409_n81), .A2(
        dp_cluster_2_mult_485_C409_n80), .A3(dp_cluster_2_mult_485_C409_n52), 
        .Z(n2639) );
  FA1D0 U1369 ( .A(dp_cluster_1_mult_513_C418_n236), .B(
        dp_cluster_1_mult_513_C418_n239), .CI(dp_cluster_1_mult_513_C418_n74), 
        .CO(dp_cluster_1_mult_513_C418_n73), .S(dp_cluster_1_N202) );
  FA1D0 U1370 ( .A(dp_cluster_3_mult_513_C415_n236), .B(
        dp_cluster_3_mult_513_C415_n239), .CI(dp_cluster_3_mult_513_C415_n74), 
        .CO(dp_cluster_3_mult_513_C415_n73), .S(dp_cluster_3_N146) );
  FA1D0 U1371 ( .A(dp_cluster_1_mult_512_C418_n236), .B(
        dp_cluster_1_mult_512_C418_n239), .CI(dp_cluster_1_mult_512_C418_n74), 
        .CO(dp_cluster_1_mult_512_C418_n73), .S(dp_cluster_1_N174) );
  FA1D0 U1372 ( .A(dp_cluster_3_mult_512_C415_n236), .B(
        dp_cluster_3_mult_512_C415_n239), .CI(dp_cluster_3_mult_512_C415_n74), 
        .CO(dp_cluster_3_mult_512_C415_n73), .S(dp_cluster_3_N118) );
  FA1D0 U1373 ( .A(dp_cluster_1_mult_513_C418_n233), .B(
        dp_cluster_1_mult_513_C418_n229), .CI(dp_cluster_1_mult_513_C418_n72), 
        .CO(dp_cluster_1_mult_513_C418_n71), .S(dp_cluster_1_N204) );
  FA1D0 U1374 ( .A(dp_cluster_0_mult_486_C412_n236), .B(
        dp_cluster_0_mult_486_C412_n239), .CI(dp_cluster_0_mult_486_C412_n74), 
        .CO(dp_cluster_0_mult_486_C412_n73), .S(dp_cluster_0_N90) );
  FA1D0 U1375 ( .A(dp_cluster_3_mult_513_C415_n233), .B(
        dp_cluster_3_mult_513_C415_n229), .CI(dp_cluster_3_mult_513_C415_n72), 
        .CO(dp_cluster_3_mult_513_C415_n71), .S(dp_cluster_3_N148) );
  FA1D0 U1376 ( .A(dp_cluster_2_mult_486_C409_n236), .B(
        dp_cluster_2_mult_486_C409_n239), .CI(dp_cluster_2_mult_486_C409_n74), 
        .CO(dp_cluster_2_mult_486_C409_n73), .S(dp_cluster_2_N34) );
  FA1D0 U1377 ( .A(dp_cluster_1_mult_512_C418_n233), .B(
        dp_cluster_1_mult_512_C418_n229), .CI(dp_cluster_1_mult_512_C418_n72), 
        .CO(dp_cluster_1_mult_512_C418_n71), .S(dp_cluster_1_N176) );
  FA1D0 U1378 ( .A(dp_cluster_3_mult_512_C415_n233), .B(
        dp_cluster_3_mult_512_C415_n229), .CI(dp_cluster_3_mult_512_C415_n72), 
        .CO(dp_cluster_3_mult_512_C415_n71), .S(dp_cluster_3_N120) );
  FA1D0 U1379 ( .A(dp_cluster_0_mult_486_C412_n233), .B(
        dp_cluster_0_mult_486_C412_n229), .CI(dp_cluster_0_mult_486_C412_n72), 
        .CO(dp_cluster_0_mult_486_C412_n71), .S(dp_cluster_0_N92) );
  FA1D0 U1380 ( .A(dp_cluster_2_mult_486_C409_n233), .B(
        dp_cluster_2_mult_486_C409_n229), .CI(dp_cluster_2_mult_486_C409_n72), 
        .CO(dp_cluster_2_mult_486_C409_n71), .S(dp_cluster_2_N36) );
  FA1D0 U1381 ( .A(dp_cluster_0_mult_485_C412_n224), .B(
        dp_cluster_0_mult_485_C412_n228), .CI(dp_cluster_0_mult_485_C412_n71), 
        .CO(dp_cluster_0_mult_485_C412_n70), .S(dp_cluster_0_N65) );
  FA1D0 U1382 ( .A(dp_cluster_2_mult_485_C409_n224), .B(
        dp_cluster_2_mult_485_C409_n228), .CI(dp_cluster_2_mult_485_C409_n71), 
        .CO(dp_cluster_2_mult_485_C409_n70), .S(dp_cluster_2_N9) );
  FA1D0 U1383 ( .A(dp_cluster_1_mult_513_C418_n217), .B(
        dp_cluster_1_mult_513_C418_n223), .CI(dp_cluster_1_mult_513_C418_n70), 
        .CO(dp_cluster_1_mult_513_C418_n69), .S(dp_cluster_1_N206) );
  FA1D0 U1384 ( .A(dp_cluster_0_mult_485_C412_n217), .B(
        dp_cluster_0_mult_485_C412_n223), .CI(dp_cluster_0_mult_485_C412_n70), 
        .CO(dp_cluster_0_mult_485_C412_n69), .S(dp_cluster_0_N66) );
  FA1D0 U1385 ( .A(dp_cluster_3_mult_513_C415_n217), .B(
        dp_cluster_3_mult_513_C415_n223), .CI(dp_cluster_3_mult_513_C415_n70), 
        .CO(dp_cluster_3_mult_513_C415_n69), .S(dp_cluster_3_N150) );
  FA1D0 U1386 ( .A(dp_cluster_2_mult_485_C409_n217), .B(
        dp_cluster_2_mult_485_C409_n223), .CI(dp_cluster_2_mult_485_C409_n70), 
        .CO(dp_cluster_2_mult_485_C409_n69), .S(dp_cluster_2_N10) );
  FA1D0 U1387 ( .A(dp_cluster_1_mult_513_C418_n211), .B(
        dp_cluster_1_mult_513_C418_n216), .CI(dp_cluster_1_mult_513_C418_n69), 
        .CO(dp_cluster_1_mult_513_C418_n68), .S(dp_cluster_1_N207) );
  FA1D0 U1388 ( .A(dp_cluster_0_mult_485_C412_n211), .B(
        dp_cluster_0_mult_485_C412_n216), .CI(dp_cluster_0_mult_485_C412_n69), 
        .CO(dp_cluster_0_mult_485_C412_n68), .S(dp_cluster_0_N67) );
  FA1D0 U1389 ( .A(dp_cluster_3_mult_513_C415_n211), .B(
        dp_cluster_3_mult_513_C415_n216), .CI(dp_cluster_3_mult_513_C415_n69), 
        .CO(dp_cluster_3_mult_513_C415_n68), .S(dp_cluster_3_N151) );
  FA1D0 U1390 ( .A(dp_cluster_2_mult_485_C409_n211), .B(
        dp_cluster_2_mult_485_C409_n216), .CI(dp_cluster_2_mult_485_C409_n69), 
        .CO(dp_cluster_2_mult_485_C409_n68), .S(dp_cluster_2_N11) );
  FA1D0 U1391 ( .A(dp_cluster_1_mult_513_C418_n203), .B(
        dp_cluster_1_mult_513_C418_n210), .CI(dp_cluster_1_mult_513_C418_n68), 
        .CO(dp_cluster_1_mult_513_C418_n67), .S(dp_cluster_1_N208) );
  FA1D0 U1392 ( .A(dp_cluster_0_mult_485_C412_n203), .B(
        dp_cluster_0_mult_485_C412_n210), .CI(dp_cluster_0_mult_485_C412_n68), 
        .CO(dp_cluster_0_mult_485_C412_n67), .S(dp_cluster_0_N68) );
  FA1D0 U1393 ( .A(dp_cluster_3_mult_513_C415_n203), .B(
        dp_cluster_3_mult_513_C415_n210), .CI(dp_cluster_3_mult_513_C415_n68), 
        .CO(dp_cluster_3_mult_513_C415_n67), .S(dp_cluster_3_N152) );
  FA1D0 U1394 ( .A(dp_cluster_2_mult_485_C409_n203), .B(
        dp_cluster_2_mult_485_C409_n210), .CI(dp_cluster_2_mult_485_C409_n68), 
        .CO(dp_cluster_2_mult_485_C409_n67), .S(dp_cluster_2_N12) );
  FA1D0 U1395 ( .A(dp_cluster_1_mult_512_C418_n195), .B(
        dp_cluster_1_mult_512_C418_n202), .CI(dp_cluster_1_mult_512_C418_n67), 
        .CO(dp_cluster_1_mult_512_C418_n66), .S(dp_cluster_1_N181) );
  FA1D0 U1396 ( .A(dp_cluster_1_mult_513_C418_n195), .B(
        dp_cluster_1_mult_513_C418_n202), .CI(dp_cluster_1_mult_513_C418_n67), 
        .CO(dp_cluster_1_mult_513_C418_n66), .S(dp_cluster_1_N209) );
  FA1D0 U1397 ( .A(dp_cluster_0_mult_485_C412_n195), .B(
        dp_cluster_0_mult_485_C412_n202), .CI(dp_cluster_0_mult_485_C412_n67), 
        .CO(dp_cluster_0_mult_485_C412_n66), .S(dp_cluster_0_N69) );
  FA1D0 U1398 ( .A(dp_cluster_3_mult_512_C415_n195), .B(
        dp_cluster_3_mult_512_C415_n202), .CI(dp_cluster_3_mult_512_C415_n67), 
        .CO(dp_cluster_3_mult_512_C415_n66), .S(dp_cluster_3_N125) );
  FA1D0 U1399 ( .A(dp_cluster_3_mult_513_C415_n195), .B(
        dp_cluster_3_mult_513_C415_n202), .CI(dp_cluster_3_mult_513_C415_n67), 
        .CO(dp_cluster_3_mult_513_C415_n66), .S(dp_cluster_3_N153) );
  FA1D0 U1400 ( .A(dp_cluster_2_mult_485_C409_n195), .B(
        dp_cluster_2_mult_485_C409_n202), .CI(dp_cluster_2_mult_485_C409_n67), 
        .CO(dp_cluster_2_mult_485_C409_n66), .S(dp_cluster_2_N13) );
  FA1D0 U1401 ( .A(dp_cluster_1_mult_513_C418_n234), .B(
        dp_cluster_1_mult_513_C418_n235), .CI(dp_cluster_1_mult_513_C418_n73), 
        .CO(dp_cluster_1_mult_513_C418_n72), .S(dp_cluster_1_N203) );
  FA1D0 U1402 ( .A(dp_cluster_3_mult_513_C415_n234), .B(
        dp_cluster_3_mult_513_C415_n235), .CI(dp_cluster_3_mult_513_C415_n73), 
        .CO(dp_cluster_3_mult_513_C415_n72), .S(dp_cluster_3_N147) );
  FA1D0 U1403 ( .A(dp_cluster_1_mult_512_C418_n234), .B(
        dp_cluster_1_mult_512_C418_n235), .CI(dp_cluster_1_mult_512_C418_n73), 
        .CO(dp_cluster_1_mult_512_C418_n72), .S(dp_cluster_1_N175) );
  FA1D0 U1404 ( .A(dp_cluster_3_mult_512_C415_n234), .B(
        dp_cluster_3_mult_512_C415_n235), .CI(dp_cluster_3_mult_512_C415_n73), 
        .CO(dp_cluster_3_mult_512_C415_n72), .S(dp_cluster_3_N119) );
  FA1D0 U1405 ( .A(dp_cluster_1_mult_513_C418_n224), .B(
        dp_cluster_1_mult_513_C418_n228), .CI(dp_cluster_1_mult_513_C418_n71), 
        .CO(dp_cluster_1_mult_513_C418_n70), .S(dp_cluster_1_N205) );
  FA1D0 U1406 ( .A(dp_cluster_3_mult_513_C415_n224), .B(
        dp_cluster_3_mult_513_C415_n228), .CI(dp_cluster_3_mult_513_C415_n71), 
        .CO(dp_cluster_3_mult_513_C415_n70), .S(dp_cluster_3_N149) );
  FA1D0 U1407 ( .A(dp_cluster_1_mult_512_C418_n224), .B(
        dp_cluster_1_mult_512_C418_n228), .CI(dp_cluster_1_mult_512_C418_n71), 
        .CO(dp_cluster_1_mult_512_C418_n70), .S(dp_cluster_1_N177) );
  FA1D0 U1408 ( .A(dp_cluster_0_mult_486_C412_n224), .B(
        dp_cluster_0_mult_486_C412_n228), .CI(dp_cluster_0_mult_486_C412_n71), 
        .CO(dp_cluster_0_mult_486_C412_n70), .S(dp_cluster_0_N93) );
  FA1D0 U1409 ( .A(dp_cluster_3_mult_512_C415_n224), .B(
        dp_cluster_3_mult_512_C415_n228), .CI(dp_cluster_3_mult_512_C415_n71), 
        .CO(dp_cluster_3_mult_512_C415_n70), .S(dp_cluster_3_N121) );
  FA1D0 U1410 ( .A(dp_cluster_2_mult_486_C409_n224), .B(
        dp_cluster_2_mult_486_C409_n228), .CI(dp_cluster_2_mult_486_C409_n71), 
        .CO(dp_cluster_2_mult_486_C409_n70), .S(dp_cluster_2_N37) );
  FA1D0 U1411 ( .A(dp_cluster_1_mult_512_C418_n217), .B(
        dp_cluster_1_mult_512_C418_n223), .CI(dp_cluster_1_mult_512_C418_n70), 
        .CO(dp_cluster_1_mult_512_C418_n69), .S(dp_cluster_1_N178) );
  FA1D0 U1412 ( .A(dp_cluster_0_mult_486_C412_n217), .B(
        dp_cluster_0_mult_486_C412_n223), .CI(dp_cluster_0_mult_486_C412_n70), 
        .CO(dp_cluster_0_mult_486_C412_n69), .S(dp_cluster_0_N94) );
  FA1D0 U1413 ( .A(dp_cluster_3_mult_512_C415_n217), .B(
        dp_cluster_3_mult_512_C415_n223), .CI(dp_cluster_3_mult_512_C415_n70), 
        .CO(dp_cluster_3_mult_512_C415_n69), .S(dp_cluster_3_N122) );
  FA1D0 U1414 ( .A(dp_cluster_2_mult_486_C409_n217), .B(
        dp_cluster_2_mult_486_C409_n223), .CI(dp_cluster_2_mult_486_C409_n70), 
        .CO(dp_cluster_2_mult_486_C409_n69), .S(dp_cluster_2_N38) );
  FA1D0 U1415 ( .A(dp_cluster_1_mult_512_C418_n211), .B(
        dp_cluster_1_mult_512_C418_n216), .CI(dp_cluster_1_mult_512_C418_n69), 
        .CO(dp_cluster_1_mult_512_C418_n68), .S(dp_cluster_1_N179) );
  FA1D0 U1416 ( .A(dp_cluster_0_mult_486_C412_n211), .B(
        dp_cluster_0_mult_486_C412_n216), .CI(dp_cluster_0_mult_486_C412_n69), 
        .CO(dp_cluster_0_mult_486_C412_n68), .S(dp_cluster_0_N95) );
  FA1D0 U1417 ( .A(dp_cluster_3_mult_512_C415_n211), .B(
        dp_cluster_3_mult_512_C415_n216), .CI(dp_cluster_3_mult_512_C415_n69), 
        .CO(dp_cluster_3_mult_512_C415_n68), .S(dp_cluster_3_N123) );
  FA1D0 U1418 ( .A(dp_cluster_2_mult_486_C409_n211), .B(
        dp_cluster_2_mult_486_C409_n216), .CI(dp_cluster_2_mult_486_C409_n69), 
        .CO(dp_cluster_2_mult_486_C409_n68), .S(dp_cluster_2_N39) );
  FA1D0 U1419 ( .A(dp_cluster_1_mult_512_C418_n203), .B(
        dp_cluster_1_mult_512_C418_n210), .CI(dp_cluster_1_mult_512_C418_n68), 
        .CO(dp_cluster_1_mult_512_C418_n67), .S(dp_cluster_1_N180) );
  FA1D0 U1420 ( .A(dp_cluster_0_mult_486_C412_n203), .B(
        dp_cluster_0_mult_486_C412_n210), .CI(dp_cluster_0_mult_486_C412_n68), 
        .CO(dp_cluster_0_mult_486_C412_n67), .S(dp_cluster_0_N96) );
  FA1D0 U1421 ( .A(dp_cluster_3_mult_512_C415_n203), .B(
        dp_cluster_3_mult_512_C415_n210), .CI(dp_cluster_3_mult_512_C415_n68), 
        .CO(dp_cluster_3_mult_512_C415_n67), .S(dp_cluster_3_N124) );
  FA1D0 U1422 ( .A(dp_cluster_2_mult_486_C409_n203), .B(
        dp_cluster_2_mult_486_C409_n210), .CI(dp_cluster_2_mult_486_C409_n68), 
        .CO(dp_cluster_2_mult_486_C409_n67), .S(dp_cluster_2_N40) );
  FA1D0 U1423 ( .A(dp_cluster_0_mult_486_C412_n195), .B(
        dp_cluster_0_mult_486_C412_n202), .CI(dp_cluster_0_mult_486_C412_n67), 
        .CO(dp_cluster_0_mult_486_C412_n66), .S(dp_cluster_0_N97) );
  FA1D0 U1424 ( .A(dp_cluster_2_mult_486_C409_n195), .B(
        dp_cluster_2_mult_486_C409_n202), .CI(dp_cluster_2_mult_486_C409_n67), 
        .CO(dp_cluster_2_mult_486_C409_n66), .S(dp_cluster_2_N41) );
  FA1D0 U1425 ( .A(dp_cluster_0_mult_485_C412_n325), .B(
        dp_cluster_0_mult_485_C412_n339), .CI(dp_cluster_0_mult_485_C412_n353), 
        .CO(dp_cluster_0_mult_485_C412_n218), .S(
        dp_cluster_0_mult_485_C412_n219) );
  OAI22D1 U1426 ( .A1(n1946), .A2(n961), .B1(n1954), .B2(n1945), .ZN(
        dp_cluster_0_mult_485_C412_n353) );
  OAI22D1 U1427 ( .A1(n1930), .A2(n960), .B1(n1936), .B2(n1929), .ZN(
        dp_cluster_0_mult_485_C412_n339) );
  OAI22D1 U1428 ( .A1(n1914), .A2(n962), .B1(n1918), .B2(n1913), .ZN(
        dp_cluster_0_mult_485_C412_n325) );
  FA1D0 U1429 ( .A(dp_cluster_2_mult_485_C409_n325), .B(
        dp_cluster_2_mult_485_C409_n339), .CI(dp_cluster_2_mult_485_C409_n353), 
        .CO(dp_cluster_2_mult_485_C409_n218), .S(
        dp_cluster_2_mult_485_C409_n219) );
  OAI22D1 U1430 ( .A1(n2597), .A2(n985), .B1(n2605), .B2(n2596), .ZN(
        dp_cluster_2_mult_485_C409_n353) );
  OAI22D1 U1431 ( .A1(n2581), .A2(n984), .B1(n2587), .B2(n2580), .ZN(
        dp_cluster_2_mult_485_C409_n339) );
  OAI22D1 U1432 ( .A1(n2565), .A2(n986), .B1(n2569), .B2(n2564), .ZN(
        dp_cluster_2_mult_485_C409_n325) );
  FA1D0 U1433 ( .A(dp_cluster_0_mult_486_C412_n325), .B(
        dp_cluster_0_mult_486_C412_n339), .CI(dp_cluster_0_mult_486_C412_n353), 
        .CO(dp_cluster_0_mult_486_C412_n218), .S(
        dp_cluster_0_mult_486_C412_n219) );
  OAI22D1 U1434 ( .A1(n1794), .A2(n955), .B1(n1802), .B2(n1793), .ZN(
        dp_cluster_0_mult_486_C412_n353) );
  OAI22D1 U1435 ( .A1(n1778), .A2(n954), .B1(n1784), .B2(n1777), .ZN(
        dp_cluster_0_mult_486_C412_n339) );
  OAI22D1 U1436 ( .A1(n1762), .A2(n956), .B1(n1766), .B2(n1761), .ZN(
        dp_cluster_0_mult_486_C412_n325) );
  FA1D0 U1437 ( .A(dp_cluster_2_mult_486_C409_n325), .B(
        dp_cluster_2_mult_486_C409_n339), .CI(dp_cluster_2_mult_486_C409_n353), 
        .CO(dp_cluster_2_mult_486_C409_n218), .S(
        dp_cluster_2_mult_486_C409_n219) );
  OAI22D1 U1438 ( .A1(n2445), .A2(n979), .B1(n2453), .B2(n2444), .ZN(
        dp_cluster_2_mult_486_C409_n353) );
  OAI22D1 U1439 ( .A1(n2429), .A2(n978), .B1(n2435), .B2(n2428), .ZN(
        dp_cluster_2_mult_486_C409_n339) );
  OAI22D1 U1440 ( .A1(n2413), .A2(n980), .B1(n2417), .B2(n2412), .ZN(
        dp_cluster_2_mult_486_C409_n325) );
  CKBD1 U1441 ( .I(n1305), .Z(n1086) );
  CKBD1 U1442 ( .I(n1272), .Z(n1064) );
  CKBD1 U1443 ( .I(n1175), .Z(n1042) );
  CKBD1 U1444 ( .I(n1136), .Z(n1020) );
  OAI22D1 U1445 ( .A1(n2229), .A2(n974), .B1(n2244), .B2(n2228), .ZN(
        dp_cluster_1_mult_512_C418_n314) );
  OAI22D1 U1446 ( .A1(n2215), .A2(n976), .B1(n2304), .B2(n2214), .ZN(
        dp_cluster_1_mult_512_C418_n299) );
  OAI22D1 U1447 ( .A1(n2203), .A2(n971), .B1(n2300), .B2(n2202), .ZN(
        dp_cluster_1_mult_512_C418_n285) );
  OAI22D1 U1448 ( .A1(n2077), .A2(n968), .B1(n2092), .B2(n2076), .ZN(
        dp_cluster_1_mult_513_C418_n314) );
  OAI22D1 U1449 ( .A1(n2063), .A2(n970), .B1(n2152), .B2(n2062), .ZN(
        dp_cluster_1_mult_513_C418_n299) );
  OAI22D1 U1450 ( .A1(n2051), .A2(n965), .B1(n2148), .B2(n2050), .ZN(
        dp_cluster_1_mult_513_C418_n285) );
  OAI22D1 U1451 ( .A1(n1751), .A2(n956), .B1(n1766), .B2(n1750), .ZN(
        dp_cluster_0_mult_486_C412_n314) );
  OAI22D1 U1452 ( .A1(n1737), .A2(n958), .B1(n1826), .B2(n1736), .ZN(
        dp_cluster_0_mult_486_C412_n299) );
  OAI22D1 U1453 ( .A1(n1725), .A2(n953), .B1(n1822), .B2(n1724), .ZN(
        dp_cluster_0_mult_486_C412_n285) );
  OAI22D1 U1454 ( .A1(n1903), .A2(n962), .B1(n1918), .B2(n1902), .ZN(
        dp_cluster_0_mult_485_C412_n314) );
  OAI22D1 U1455 ( .A1(n1889), .A2(n964), .B1(n1978), .B2(n1888), .ZN(
        dp_cluster_0_mult_485_C412_n299) );
  OAI22D1 U1456 ( .A1(n1877), .A2(n959), .B1(n1974), .B2(n1876), .ZN(
        dp_cluster_0_mult_485_C412_n285) );
  OAI22D1 U1457 ( .A1(n2880), .A2(n998), .B1(n2895), .B2(n2879), .ZN(
        dp_cluster_3_mult_512_C415_n314) );
  OAI22D1 U1458 ( .A1(n2866), .A2(n1000), .B1(n2955), .B2(n2865), .ZN(
        dp_cluster_3_mult_512_C415_n299) );
  OAI22D1 U1459 ( .A1(n2854), .A2(n995), .B1(n2951), .B2(n2853), .ZN(
        dp_cluster_3_mult_512_C415_n285) );
  OAI22D1 U1460 ( .A1(n2728), .A2(n992), .B1(n2743), .B2(n2727), .ZN(
        dp_cluster_3_mult_513_C415_n314) );
  OAI22D1 U1461 ( .A1(n2714), .A2(n994), .B1(n2803), .B2(n2713), .ZN(
        dp_cluster_3_mult_513_C415_n299) );
  OAI22D1 U1462 ( .A1(n2702), .A2(n989), .B1(n2799), .B2(n2701), .ZN(
        dp_cluster_3_mult_513_C415_n285) );
  OAI22D1 U1463 ( .A1(n2402), .A2(n980), .B1(n2417), .B2(n2401), .ZN(
        dp_cluster_2_mult_486_C409_n314) );
  OAI22D1 U1464 ( .A1(n2388), .A2(n982), .B1(n2477), .B2(n2387), .ZN(
        dp_cluster_2_mult_486_C409_n299) );
  OAI22D1 U1465 ( .A1(n2376), .A2(n977), .B1(n2473), .B2(n2375), .ZN(
        dp_cluster_2_mult_486_C409_n285) );
  OAI22D1 U1466 ( .A1(n2554), .A2(n986), .B1(n2569), .B2(n2553), .ZN(
        dp_cluster_2_mult_485_C409_n314) );
  OAI22D1 U1467 ( .A1(n2540), .A2(n988), .B1(n2629), .B2(n2539), .ZN(
        dp_cluster_2_mult_485_C409_n299) );
  OAI22D1 U1468 ( .A1(n2528), .A2(n983), .B1(n2625), .B2(n2527), .ZN(
        dp_cluster_2_mult_485_C409_n285) );
  FA1D0 U1469 ( .A(dp_cluster_0_mult_485_C412_n236), .B(
        dp_cluster_0_mult_485_C412_n239), .CI(dp_cluster_0_mult_485_C412_n74), 
        .CO(dp_cluster_0_mult_485_C412_n73), .S(dp_cluster_0_N62) );
  FA1D0 U1470 ( .A(dp_cluster_2_mult_485_C409_n236), .B(
        dp_cluster_2_mult_485_C409_n239), .CI(dp_cluster_2_mult_485_C409_n74), 
        .CO(dp_cluster_2_mult_485_C409_n73), .S(dp_cluster_2_N6) );
  FA1D0 U1471 ( .A(dp_cluster_0_mult_485_C412_n233), .B(
        dp_cluster_0_mult_485_C412_n229), .CI(dp_cluster_0_mult_485_C412_n72), 
        .CO(dp_cluster_0_mult_485_C412_n71), .S(dp_cluster_0_N64) );
  FA1D0 U1472 ( .A(dp_cluster_2_mult_485_C409_n233), .B(
        dp_cluster_2_mult_485_C409_n229), .CI(dp_cluster_2_mult_485_C409_n72), 
        .CO(dp_cluster_2_mult_485_C409_n71), .S(dp_cluster_2_N8) );
  IOA21D1 U1473 ( .A1(n2324), .A2(dp_cluster_1_N174), .B(n2323), .ZN(n2326) );
  OAI21D1 U1474 ( .A1(dp_cluster_1_N174), .A2(n2324), .B(dp_cluster_1_N202), 
        .ZN(n2323) );
  IOA21D1 U1475 ( .A1(n2322), .A2(dp_cluster_1_N173), .B(n2321), .ZN(n2324) );
  OAI21D1 U1476 ( .A1(dp_cluster_1_N173), .A2(n2322), .B(dp_cluster_1_N201), 
        .ZN(n2321) );
  IOA21D1 U1477 ( .A1(n2975), .A2(dp_cluster_3_N118), .B(n2974), .ZN(n2977) );
  OAI21D1 U1478 ( .A1(dp_cluster_3_N118), .A2(n2975), .B(dp_cluster_3_N146), 
        .ZN(n2974) );
  IOA21D1 U1479 ( .A1(n2973), .A2(dp_cluster_3_N117), .B(n2972), .ZN(n2975) );
  OAI21D1 U1480 ( .A1(dp_cluster_3_N117), .A2(n2973), .B(dp_cluster_3_N145), 
        .ZN(n2972) );
  CKBD1 U1481 ( .I(n1173), .Z(n1039) );
  CKBD1 U1482 ( .I(n1134), .Z(n1017) );
  CKBD1 U1483 ( .I(n1304), .Z(n1083) );
  CKBD1 U1484 ( .I(n1271), .Z(n1061) );
  CKBD1 U1485 ( .I(n1163), .Z(n1030) );
  CKBD1 U1486 ( .I(n1124), .Z(n1008) );
  CKBD1 U1487 ( .I(n1298), .Z(n1077) );
  CKBD1 U1488 ( .I(n1265), .Z(n1055) );
  CKBD1 U1489 ( .I(n1165), .Z(n1033) );
  CKBD1 U1490 ( .I(n1126), .Z(n1011) );
  CKBD1 U1491 ( .I(n1297), .Z(n1074) );
  CKBD1 U1492 ( .I(n1264), .Z(n1052) );
  CKBD1 U1493 ( .I(n1153), .Z(n1025) );
  CKBD1 U1494 ( .I(n1288), .Z(n1069) );
  CKBD1 U1495 ( .I(n1114), .Z(n1003) );
  CKBD1 U1496 ( .I(n1255), .Z(n1047) );
  CKBD1 U1497 ( .I(n1304), .Z(n1084) );
  CKBD1 U1498 ( .I(n1271), .Z(n1062) );
  CKBD1 U1499 ( .I(n1165), .Z(n1034) );
  CKBD1 U1500 ( .I(n1173), .Z(n1040) );
  CKBD1 U1501 ( .I(n1126), .Z(n1012) );
  CKBD1 U1502 ( .I(n1134), .Z(n1018) );
  CKBD1 U1503 ( .I(n1163), .Z(n1031) );
  CKBD1 U1504 ( .I(n1124), .Z(n1009) );
  CKBD1 U1505 ( .I(n1297), .Z(n1075) );
  CKBD1 U1506 ( .I(n1298), .Z(n1078) );
  CKBD1 U1507 ( .I(n1264), .Z(n1053) );
  CKBD1 U1508 ( .I(n1265), .Z(n1056) );
  CKBD1 U1509 ( .I(n1153), .Z(n1026) );
  CKBD1 U1510 ( .I(n1114), .Z(n1004) );
  CKBD1 U1511 ( .I(n1288), .Z(n1070) );
  CKBD1 U1512 ( .I(n1255), .Z(n1048) );
  CKBD1 U1513 ( .I(n1301), .Z(n1081) );
  CKBD1 U1514 ( .I(n1268), .Z(n1059) );
  CKBD1 U1515 ( .I(n1169), .Z(n1037) );
  CKBD1 U1516 ( .I(n1130), .Z(n1015) );
  CKBD1 U1517 ( .I(n1169), .Z(n1036) );
  CKBD1 U1518 ( .I(n1130), .Z(n1014) );
  CKBD1 U1519 ( .I(n1301), .Z(n1080) );
  CKBD1 U1520 ( .I(n1268), .Z(n1058) );
  CKBD1 U1521 ( .I(n1159), .Z(n1028) );
  CKBD1 U1522 ( .I(n1294), .Z(n1072) );
  CKBD1 U1523 ( .I(n1120), .Z(n1006) );
  CKBD1 U1524 ( .I(n1261), .Z(n1050) );
  CKBD1 U1525 ( .I(n1175), .Z(n1043) );
  CKBD1 U1526 ( .I(n1136), .Z(n1021) );
  CKBD1 U1527 ( .I(n1305), .Z(n1087) );
  CKBD1 U1528 ( .I(n1272), .Z(n1065) );
  CKBD1 U1529 ( .I(n1285), .Z(n1067) );
  CKBD1 U1530 ( .I(n1152), .Z(n1023) );
  CKBD1 U1531 ( .I(n1252), .Z(n1045) );
  CKBD1 U1532 ( .I(n1113), .Z(n1001) );
  CKBD1 U1533 ( .I(n1294), .Z(n1073) );
  CKBD1 U1534 ( .I(n1159), .Z(n1029) );
  CKBD1 U1535 ( .I(n1261), .Z(n1051) );
  CKBD1 U1536 ( .I(n1120), .Z(n1007) );
  FA1D0 U1537 ( .A(dp_cluster_1_mult_512_C418_n269), .B(
        dp_cluster_1_mult_512_C418_n255), .CI(n1162), .CO(
        dp_cluster_1_mult_512_C418_n96), .S(dp_cluster_1_mult_512_C418_n97) );
  INVD1 U1538 ( .I(dp_cluster_1_mult_512_C418_n98), .ZN(n1162) );
  OAI22D1 U1539 ( .A1(n2188), .A2(n975), .B1(n2310), .B2(n2187), .ZN(
        dp_cluster_1_mult_512_C418_n269) );
  OAI22D1 U1540 ( .A1(n2176), .A2(n2306), .B1(n2307), .B2(n2175), .ZN(
        dp_cluster_1_mult_512_C418_n255) );
  FA1D0 U1541 ( .A(dp_cluster_1_mult_513_C418_n269), .B(
        dp_cluster_1_mult_513_C418_n255), .CI(n1296), .CO(
        dp_cluster_1_mult_513_C418_n96), .S(dp_cluster_1_mult_513_C418_n97) );
  INVD1 U1542 ( .I(dp_cluster_1_mult_513_C418_n98), .ZN(n1296) );
  OAI22D1 U1543 ( .A1(n2036), .A2(n969), .B1(n2158), .B2(n2035), .ZN(
        dp_cluster_1_mult_513_C418_n269) );
  OAI22D1 U1544 ( .A1(n2024), .A2(n2154), .B1(n2155), .B2(n2023), .ZN(
        dp_cluster_1_mult_513_C418_n255) );
  FA1D0 U1545 ( .A(dp_cluster_0_mult_486_C412_n269), .B(
        dp_cluster_0_mult_486_C412_n255), .CI(n1295), .CO(
        dp_cluster_0_mult_486_C412_n96), .S(dp_cluster_0_mult_486_C412_n97) );
  INVD1 U1546 ( .I(dp_cluster_0_mult_486_C412_n98), .ZN(n1295) );
  OAI22D1 U1547 ( .A1(n1710), .A2(n957), .B1(n1832), .B2(n1709), .ZN(
        dp_cluster_0_mult_486_C412_n269) );
  OAI22D1 U1548 ( .A1(n1698), .A2(n1828), .B1(n1829), .B2(n1697), .ZN(
        dp_cluster_0_mult_486_C412_n255) );
  FA1D0 U1549 ( .A(dp_cluster_0_mult_485_C412_n269), .B(
        dp_cluster_0_mult_485_C412_n255), .CI(n1161), .CO(
        dp_cluster_0_mult_485_C412_n96), .S(dp_cluster_0_mult_485_C412_n97) );
  INVD1 U1550 ( .I(dp_cluster_0_mult_485_C412_n98), .ZN(n1161) );
  OAI22D1 U1551 ( .A1(n1862), .A2(n963), .B1(n1984), .B2(n1861), .ZN(
        dp_cluster_0_mult_485_C412_n269) );
  OAI22D1 U1552 ( .A1(n1850), .A2(n1980), .B1(n1981), .B2(n1849), .ZN(
        dp_cluster_0_mult_485_C412_n255) );
  FA1D0 U1553 ( .A(dp_cluster_3_mult_512_C415_n269), .B(
        dp_cluster_3_mult_512_C415_n255), .CI(n1123), .CO(
        dp_cluster_3_mult_512_C415_n96), .S(dp_cluster_3_mult_512_C415_n97) );
  INVD1 U1554 ( .I(dp_cluster_3_mult_512_C415_n98), .ZN(n1123) );
  OAI22D1 U1555 ( .A1(n2839), .A2(n999), .B1(n2961), .B2(n2838), .ZN(
        dp_cluster_3_mult_512_C415_n269) );
  OAI22D1 U1556 ( .A1(n2827), .A2(n2957), .B1(n2958), .B2(n2826), .ZN(
        dp_cluster_3_mult_512_C415_n255) );
  FA1D0 U1557 ( .A(dp_cluster_3_mult_513_C415_n269), .B(
        dp_cluster_3_mult_513_C415_n255), .CI(n1263), .CO(
        dp_cluster_3_mult_513_C415_n96), .S(dp_cluster_3_mult_513_C415_n97) );
  INVD1 U1558 ( .I(dp_cluster_3_mult_513_C415_n98), .ZN(n1263) );
  OAI22D1 U1559 ( .A1(n2687), .A2(n993), .B1(n2809), .B2(n2686), .ZN(
        dp_cluster_3_mult_513_C415_n269) );
  OAI22D1 U1560 ( .A1(n2675), .A2(n2805), .B1(n2806), .B2(n2674), .ZN(
        dp_cluster_3_mult_513_C415_n255) );
  FA1D0 U1561 ( .A(dp_cluster_2_mult_486_C409_n269), .B(
        dp_cluster_2_mult_486_C409_n255), .CI(n1262), .CO(
        dp_cluster_2_mult_486_C409_n96), .S(dp_cluster_2_mult_486_C409_n97) );
  INVD1 U1562 ( .I(dp_cluster_2_mult_486_C409_n98), .ZN(n1262) );
  OAI22D1 U1563 ( .A1(n2361), .A2(n981), .B1(n2483), .B2(n2360), .ZN(
        dp_cluster_2_mult_486_C409_n269) );
  OAI22D1 U1564 ( .A1(n2349), .A2(n2479), .B1(n2480), .B2(n2348), .ZN(
        dp_cluster_2_mult_486_C409_n255) );
  FA1D0 U1565 ( .A(dp_cluster_2_mult_485_C409_n269), .B(
        dp_cluster_2_mult_485_C409_n255), .CI(n1122), .CO(
        dp_cluster_2_mult_485_C409_n96), .S(dp_cluster_2_mult_485_C409_n97) );
  INVD1 U1566 ( .I(dp_cluster_2_mult_485_C409_n98), .ZN(n1122) );
  OAI22D1 U1567 ( .A1(n2513), .A2(n987), .B1(n2635), .B2(n2512), .ZN(
        dp_cluster_2_mult_485_C409_n269) );
  OAI22D1 U1568 ( .A1(n2501), .A2(n2631), .B1(n2632), .B2(n2500), .ZN(
        dp_cluster_2_mult_485_C409_n255) );
  FA1D0 U1569 ( .A(dp_cluster_0_mult_486_C412_n84), .B(
        dp_cluster_0_mult_486_C412_n82), .CI(dp_cluster_0_mult_486_C412_n53), 
        .CO(dp_cluster_0_mult_486_C412_n52), .S(dp_cluster_0_N111) );
  FA1D0 U1570 ( .A(dp_cluster_2_mult_486_C409_n84), .B(
        dp_cluster_2_mult_486_C409_n82), .CI(dp_cluster_2_mult_486_C409_n53), 
        .CO(dp_cluster_2_mult_486_C409_n52), .S(dp_cluster_2_N55) );
  FA1D0 U1571 ( .A(dp_cluster_1_mult_512_C418_n84), .B(
        dp_cluster_1_mult_512_C418_n82), .CI(dp_cluster_1_mult_512_C418_n53), 
        .CO(dp_cluster_1_mult_512_C418_n52), .S(dp_cluster_1_N195) );
  FA1D0 U1572 ( .A(dp_cluster_1_mult_513_C418_n84), .B(
        dp_cluster_1_mult_513_C418_n82), .CI(dp_cluster_1_mult_513_C418_n53), 
        .CO(dp_cluster_1_mult_513_C418_n52), .S(dp_cluster_1_N223) );
  FA1D0 U1573 ( .A(dp_cluster_0_mult_485_C412_n84), .B(
        dp_cluster_0_mult_485_C412_n82), .CI(dp_cluster_0_mult_485_C412_n53), 
        .CO(dp_cluster_0_mult_485_C412_n52), .S(dp_cluster_0_N83) );
  FA1D0 U1574 ( .A(dp_cluster_3_mult_512_C415_n84), .B(
        dp_cluster_3_mult_512_C415_n82), .CI(dp_cluster_3_mult_512_C415_n53), 
        .CO(dp_cluster_3_mult_512_C415_n52), .S(dp_cluster_3_N139) );
  FA1D0 U1575 ( .A(dp_cluster_3_mult_513_C415_n84), .B(
        dp_cluster_3_mult_513_C415_n82), .CI(dp_cluster_3_mult_513_C415_n53), 
        .CO(dp_cluster_3_mult_513_C415_n52), .S(dp_cluster_3_N167) );
  FA1D0 U1576 ( .A(dp_cluster_2_mult_485_C409_n84), .B(
        dp_cluster_2_mult_485_C409_n82), .CI(dp_cluster_2_mult_485_C409_n53), 
        .CO(dp_cluster_2_mult_485_C409_n52), .S(dp_cluster_2_N27) );
  FA1D0 U1577 ( .A(dp_cluster_1_mult_512_C418_n315), .B(
        dp_cluster_1_mult_512_C418_n273), .CI(n1168), .CO(
        dp_cluster_1_mult_512_C418_n128), .S(dp_cluster_1_mult_512_C418_n129)
         );
  INVD1 U1578 ( .I(dp_cluster_1_mult_512_C418_n130), .ZN(n1168) );
  OAI22D1 U1579 ( .A1(n2230), .A2(n974), .B1(n2244), .B2(n2229), .ZN(
        dp_cluster_1_mult_512_C418_n315) );
  OAI22D1 U1580 ( .A1(n2192), .A2(n975), .B1(n2310), .B2(n2191), .ZN(
        dp_cluster_1_mult_512_C418_n273) );
  FA1D0 U1581 ( .A(dp_cluster_1_mult_513_C418_n315), .B(
        dp_cluster_1_mult_513_C418_n273), .CI(n1300), .CO(
        dp_cluster_1_mult_513_C418_n128), .S(dp_cluster_1_mult_513_C418_n129)
         );
  INVD1 U1582 ( .I(dp_cluster_1_mult_513_C418_n130), .ZN(n1300) );
  OAI22D1 U1583 ( .A1(n2078), .A2(n968), .B1(n2092), .B2(n2077), .ZN(
        dp_cluster_1_mult_513_C418_n315) );
  OAI22D1 U1584 ( .A1(n2040), .A2(n969), .B1(n2158), .B2(n2039), .ZN(
        dp_cluster_1_mult_513_C418_n273) );
  FA1D0 U1585 ( .A(dp_cluster_0_mult_486_C412_n315), .B(
        dp_cluster_0_mult_486_C412_n273), .CI(n1299), .CO(
        dp_cluster_0_mult_486_C412_n128), .S(dp_cluster_0_mult_486_C412_n129)
         );
  INVD1 U1586 ( .I(dp_cluster_0_mult_486_C412_n130), .ZN(n1299) );
  OAI22D1 U1587 ( .A1(n1752), .A2(n956), .B1(n1766), .B2(n1751), .ZN(
        dp_cluster_0_mult_486_C412_n315) );
  OAI22D1 U1588 ( .A1(n1714), .A2(n957), .B1(n1832), .B2(n1713), .ZN(
        dp_cluster_0_mult_486_C412_n273) );
  FA1D0 U1589 ( .A(dp_cluster_0_mult_485_C412_n315), .B(
        dp_cluster_0_mult_485_C412_n273), .CI(n1166), .CO(
        dp_cluster_0_mult_485_C412_n128), .S(dp_cluster_0_mult_485_C412_n129)
         );
  INVD1 U1590 ( .I(dp_cluster_0_mult_485_C412_n130), .ZN(n1166) );
  OAI22D1 U1591 ( .A1(n1904), .A2(n962), .B1(n1918), .B2(n1903), .ZN(
        dp_cluster_0_mult_485_C412_n315) );
  OAI22D1 U1592 ( .A1(n1866), .A2(n963), .B1(n1984), .B2(n1865), .ZN(
        dp_cluster_0_mult_485_C412_n273) );
  FA1D0 U1593 ( .A(dp_cluster_3_mult_512_C415_n315), .B(
        dp_cluster_3_mult_512_C415_n273), .CI(n1129), .CO(
        dp_cluster_3_mult_512_C415_n128), .S(dp_cluster_3_mult_512_C415_n129)
         );
  INVD1 U1594 ( .I(dp_cluster_3_mult_512_C415_n130), .ZN(n1129) );
  OAI22D1 U1595 ( .A1(n2881), .A2(n998), .B1(n2895), .B2(n2880), .ZN(
        dp_cluster_3_mult_512_C415_n315) );
  OAI22D1 U1596 ( .A1(n2843), .A2(n999), .B1(n2961), .B2(n2842), .ZN(
        dp_cluster_3_mult_512_C415_n273) );
  FA1D0 U1597 ( .A(dp_cluster_3_mult_513_C415_n315), .B(
        dp_cluster_3_mult_513_C415_n273), .CI(n1267), .CO(
        dp_cluster_3_mult_513_C415_n128), .S(dp_cluster_3_mult_513_C415_n129)
         );
  INVD1 U1598 ( .I(dp_cluster_3_mult_513_C415_n130), .ZN(n1267) );
  OAI22D1 U1599 ( .A1(n2729), .A2(n992), .B1(n2743), .B2(n2728), .ZN(
        dp_cluster_3_mult_513_C415_n315) );
  OAI22D1 U1600 ( .A1(n2691), .A2(n993), .B1(n2809), .B2(n2690), .ZN(
        dp_cluster_3_mult_513_C415_n273) );
  FA1D0 U1601 ( .A(dp_cluster_2_mult_486_C409_n315), .B(
        dp_cluster_2_mult_486_C409_n273), .CI(n1266), .CO(
        dp_cluster_2_mult_486_C409_n128), .S(dp_cluster_2_mult_486_C409_n129)
         );
  INVD1 U1602 ( .I(dp_cluster_2_mult_486_C409_n130), .ZN(n1266) );
  OAI22D1 U1603 ( .A1(n2403), .A2(n980), .B1(n2417), .B2(n2402), .ZN(
        dp_cluster_2_mult_486_C409_n315) );
  OAI22D1 U1604 ( .A1(n2365), .A2(n981), .B1(n2483), .B2(n2364), .ZN(
        dp_cluster_2_mult_486_C409_n273) );
  FA1D0 U1605 ( .A(dp_cluster_2_mult_485_C409_n315), .B(
        dp_cluster_2_mult_485_C409_n273), .CI(n1127), .CO(
        dp_cluster_2_mult_485_C409_n128), .S(dp_cluster_2_mult_485_C409_n129)
         );
  INVD1 U1606 ( .I(dp_cluster_2_mult_485_C409_n130), .ZN(n1127) );
  OAI22D1 U1607 ( .A1(n2555), .A2(n986), .B1(n2569), .B2(n2554), .ZN(
        dp_cluster_2_mult_485_C409_n315) );
  OAI22D1 U1608 ( .A1(n2517), .A2(n987), .B1(n2635), .B2(n2516), .ZN(
        dp_cluster_2_mult_485_C409_n273) );
  FA1D0 U1609 ( .A(dp_cluster_0_mult_486_C412_n234), .B(
        dp_cluster_0_mult_486_C412_n235), .CI(dp_cluster_0_mult_486_C412_n73), 
        .CO(dp_cluster_0_mult_486_C412_n72), .S(dp_cluster_0_N91) );
  FA1D0 U1610 ( .A(dp_cluster_2_mult_486_C409_n234), .B(
        dp_cluster_2_mult_486_C409_n235), .CI(dp_cluster_2_mult_486_C409_n73), 
        .CO(dp_cluster_2_mult_486_C409_n72), .S(dp_cluster_2_N35) );
  FA1D0 U1611 ( .A(dp_cluster_1_mult_513_C418_n340), .B(
        dp_cluster_1_mult_513_C418_n311), .CI(dp_cluster_1_mult_513_C418_n326), 
        .CO(dp_cluster_1_mult_513_C418_n225), .S(
        dp_cluster_1_mult_513_C418_n226) );
  OAI22D1 U1612 ( .A1(n2105), .A2(n966), .B1(n2110), .B2(n2104), .ZN(
        dp_cluster_1_mult_513_C418_n340) );
  OAI22D1 U1613 ( .A1(n2089), .A2(n968), .B1(n2092), .B2(n2088), .ZN(
        dp_cluster_1_mult_513_C418_n326) );
  NR2D1 U1614 ( .A1(n2152), .A2(n1092), .ZN(dp_cluster_1_mult_513_C418_n311)
         );
  FA1D0 U1615 ( .A(dp_cluster_0_mult_485_C412_n340), .B(
        dp_cluster_0_mult_485_C412_n311), .CI(dp_cluster_0_mult_485_C412_n326), 
        .CO(dp_cluster_0_mult_485_C412_n225), .S(
        dp_cluster_0_mult_485_C412_n226) );
  OAI22D1 U1616 ( .A1(n1931), .A2(n960), .B1(n1936), .B2(n1930), .ZN(
        dp_cluster_0_mult_485_C412_n340) );
  OAI22D1 U1617 ( .A1(n1915), .A2(n962), .B1(n1918), .B2(n1914), .ZN(
        dp_cluster_0_mult_485_C412_n326) );
  NR2D1 U1618 ( .A1(n1978), .A2(n1093), .ZN(dp_cluster_0_mult_485_C412_n311)
         );
  FA1D0 U1619 ( .A(dp_cluster_3_mult_513_C415_n340), .B(
        dp_cluster_3_mult_513_C415_n311), .CI(dp_cluster_3_mult_513_C415_n326), 
        .CO(dp_cluster_3_mult_513_C415_n225), .S(
        dp_cluster_3_mult_513_C415_n226) );
  OAI22D1 U1620 ( .A1(n2756), .A2(n990), .B1(n2761), .B2(n2755), .ZN(
        dp_cluster_3_mult_513_C415_n340) );
  OAI22D1 U1621 ( .A1(n2740), .A2(n992), .B1(n2743), .B2(n2739), .ZN(
        dp_cluster_3_mult_513_C415_n326) );
  NR2D1 U1622 ( .A1(n2803), .A2(n1089), .ZN(dp_cluster_3_mult_513_C415_n311)
         );
  FA1D0 U1623 ( .A(dp_cluster_2_mult_485_C409_n340), .B(
        dp_cluster_2_mult_485_C409_n311), .CI(dp_cluster_2_mult_485_C409_n326), 
        .CO(dp_cluster_2_mult_485_C409_n225), .S(
        dp_cluster_2_mult_485_C409_n226) );
  OAI22D1 U1624 ( .A1(n2582), .A2(n984), .B1(n2587), .B2(n2581), .ZN(
        dp_cluster_2_mult_485_C409_n340) );
  OAI22D1 U1625 ( .A1(n2566), .A2(n986), .B1(n2569), .B2(n2565), .ZN(
        dp_cluster_2_mult_485_C409_n326) );
  NR2D1 U1626 ( .A1(n2629), .A2(n1090), .ZN(dp_cluster_2_mult_485_C409_n311)
         );
  FA1D0 U1627 ( .A(dp_cluster_1_mult_512_C418_n340), .B(
        dp_cluster_1_mult_512_C418_n311), .CI(dp_cluster_1_mult_512_C418_n326), 
        .CO(dp_cluster_1_mult_512_C418_n225), .S(
        dp_cluster_1_mult_512_C418_n226) );
  OAI22D1 U1628 ( .A1(n2257), .A2(n972), .B1(n2262), .B2(n2256), .ZN(
        dp_cluster_1_mult_512_C418_n340) );
  OAI22D1 U1629 ( .A1(n2241), .A2(n974), .B1(n2244), .B2(n2240), .ZN(
        dp_cluster_1_mult_512_C418_n326) );
  NR2D1 U1630 ( .A1(n2304), .A2(n1098), .ZN(dp_cluster_1_mult_512_C418_n311)
         );
  FA1D0 U1631 ( .A(dp_cluster_0_mult_486_C412_n340), .B(
        dp_cluster_0_mult_486_C412_n311), .CI(dp_cluster_0_mult_486_C412_n326), 
        .CO(dp_cluster_0_mult_486_C412_n225), .S(
        dp_cluster_0_mult_486_C412_n226) );
  OAI22D1 U1632 ( .A1(n1779), .A2(n954), .B1(n1784), .B2(n1778), .ZN(
        dp_cluster_0_mult_486_C412_n340) );
  OAI22D1 U1633 ( .A1(n1763), .A2(n956), .B1(n1766), .B2(n1762), .ZN(
        dp_cluster_0_mult_486_C412_n326) );
  NR2D1 U1634 ( .A1(n1826), .A2(n1099), .ZN(dp_cluster_0_mult_486_C412_n311)
         );
  FA1D0 U1635 ( .A(dp_cluster_3_mult_512_C415_n340), .B(
        dp_cluster_3_mult_512_C415_n311), .CI(dp_cluster_3_mult_512_C415_n326), 
        .CO(dp_cluster_3_mult_512_C415_n225), .S(
        dp_cluster_3_mult_512_C415_n226) );
  OAI22D1 U1636 ( .A1(n2908), .A2(n996), .B1(n2913), .B2(n2907), .ZN(
        dp_cluster_3_mult_512_C415_n340) );
  OAI22D1 U1637 ( .A1(n2892), .A2(n998), .B1(n2895), .B2(n2891), .ZN(
        dp_cluster_3_mult_512_C415_n326) );
  NR2D1 U1638 ( .A1(n2955), .A2(n1095), .ZN(dp_cluster_3_mult_512_C415_n311)
         );
  FA1D0 U1639 ( .A(dp_cluster_2_mult_486_C409_n340), .B(
        dp_cluster_2_mult_486_C409_n311), .CI(dp_cluster_2_mult_486_C409_n326), 
        .CO(dp_cluster_2_mult_486_C409_n225), .S(
        dp_cluster_2_mult_486_C409_n226) );
  OAI22D1 U1640 ( .A1(n2430), .A2(n978), .B1(n2435), .B2(n2429), .ZN(
        dp_cluster_2_mult_486_C409_n340) );
  OAI22D1 U1641 ( .A1(n2414), .A2(n980), .B1(n2417), .B2(n2413), .ZN(
        dp_cluster_2_mult_486_C409_n326) );
  NR2D1 U1642 ( .A1(n2477), .A2(n1096), .ZN(dp_cluster_2_mult_486_C409_n311)
         );
  CKBD1 U1643 ( .I(n1285), .Z(n1068) );
  CKBD1 U1644 ( .I(n1152), .Z(n1024) );
  CKBD1 U1645 ( .I(n1252), .Z(n1046) );
  CKBD1 U1646 ( .I(n1113), .Z(n1002) );
  CKBD1 U1647 ( .I(n1305), .Z(n1088) );
  CKBD1 U1648 ( .I(n1175), .Z(n1044) );
  CKBD1 U1649 ( .I(n1272), .Z(n1066) );
  CKBD1 U1650 ( .I(n1136), .Z(n1022) );
  CKBD1 U1651 ( .I(n1169), .Z(n1038) );
  CKBD1 U1652 ( .I(n1130), .Z(n1016) );
  CKBD1 U1653 ( .I(n1301), .Z(n1082) );
  CKBD1 U1654 ( .I(n1268), .Z(n1060) );
  CKBD1 U1655 ( .I(n1163), .Z(n1032) );
  CKBD1 U1656 ( .I(n1124), .Z(n1010) );
  CKBD1 U1657 ( .I(n1288), .Z(n1071) );
  CKBD1 U1658 ( .I(n1153), .Z(n1027) );
  CKBD1 U1659 ( .I(n1255), .Z(n1049) );
  CKBD1 U1660 ( .I(n1114), .Z(n1005) );
  CKBD1 U1661 ( .I(n1173), .Z(n1041) );
  CKBD1 U1662 ( .I(n1134), .Z(n1019) );
  CKBD1 U1663 ( .I(n1304), .Z(n1085) );
  CKBD1 U1664 ( .I(n1271), .Z(n1063) );
  CKBD1 U1665 ( .I(n1165), .Z(n1035) );
  CKBD1 U1666 ( .I(n1298), .Z(n1079) );
  CKBD1 U1667 ( .I(n1126), .Z(n1013) );
  CKBD1 U1668 ( .I(n1265), .Z(n1057) );
  CKBD1 U1669 ( .I(n1297), .Z(n1076) );
  CKBD1 U1670 ( .I(n1264), .Z(n1054) );
  OAI22D1 U1671 ( .A1(n2199), .A2(n971), .B1(n2300), .B2(n2298), .ZN(
        dp_cluster_1_mult_512_C418_n282) );
  OAI22D1 U1672 ( .A1(n2047), .A2(n965), .B1(n2148), .B2(n2146), .ZN(
        dp_cluster_1_mult_513_C418_n282) );
  OAI22D1 U1673 ( .A1(n1721), .A2(n953), .B1(n1822), .B2(n1820), .ZN(
        dp_cluster_0_mult_486_C412_n282) );
  OAI22D1 U1674 ( .A1(n1873), .A2(n959), .B1(n1974), .B2(n1972), .ZN(
        dp_cluster_0_mult_485_C412_n282) );
  OAI22D1 U1675 ( .A1(n2850), .A2(n995), .B1(n2951), .B2(n2949), .ZN(
        dp_cluster_3_mult_512_C415_n282) );
  OAI22D1 U1676 ( .A1(n2698), .A2(n989), .B1(n2799), .B2(n2797), .ZN(
        dp_cluster_3_mult_513_C415_n282) );
  OAI22D1 U1677 ( .A1(n2372), .A2(n977), .B1(n2473), .B2(n2471), .ZN(
        dp_cluster_2_mult_486_C409_n282) );
  OAI22D1 U1678 ( .A1(n2524), .A2(n983), .B1(n2625), .B2(n2623), .ZN(
        dp_cluster_2_mult_485_C409_n282) );
  INVD1 U1679 ( .I(dp_cluster_1_mult_512_C418_n86), .ZN(n1158) );
  OAI22D1 U1680 ( .A1(n2186), .A2(n975), .B1(n2310), .B2(n2185), .ZN(
        dp_cluster_1_mult_512_C418_n267) );
  OAI22D1 U1681 ( .A1(n2174), .A2(n2306), .B1(n2307), .B2(n2173), .ZN(
        dp_cluster_1_mult_512_C418_n253) );
  INVD1 U1682 ( .I(dp_cluster_1_mult_513_C418_n86), .ZN(n1293) );
  OAI22D1 U1683 ( .A1(n2034), .A2(n969), .B1(n2158), .B2(n2033), .ZN(
        dp_cluster_1_mult_513_C418_n267) );
  OAI22D1 U1684 ( .A1(n2022), .A2(n2154), .B1(n2155), .B2(n2021), .ZN(
        dp_cluster_1_mult_513_C418_n253) );
  INVD1 U1685 ( .I(dp_cluster_0_mult_486_C412_n86), .ZN(n1291) );
  OAI22D1 U1686 ( .A1(n1708), .A2(n957), .B1(n1832), .B2(n1707), .ZN(
        dp_cluster_0_mult_486_C412_n267) );
  OAI22D1 U1687 ( .A1(n1696), .A2(n1828), .B1(n1829), .B2(n1695), .ZN(
        dp_cluster_0_mult_486_C412_n253) );
  INVD1 U1688 ( .I(dp_cluster_0_mult_485_C412_n86), .ZN(n1156) );
  OAI22D1 U1689 ( .A1(n1860), .A2(n963), .B1(n1984), .B2(n1859), .ZN(
        dp_cluster_0_mult_485_C412_n267) );
  OAI22D1 U1690 ( .A1(n1848), .A2(n1980), .B1(n1981), .B2(n1847), .ZN(
        dp_cluster_0_mult_485_C412_n253) );
  INVD1 U1691 ( .I(dp_cluster_3_mult_512_C415_n86), .ZN(n1119) );
  OAI22D1 U1692 ( .A1(n2837), .A2(n999), .B1(n2961), .B2(n2836), .ZN(
        dp_cluster_3_mult_512_C415_n267) );
  OAI22D1 U1693 ( .A1(n2825), .A2(n2957), .B1(n2958), .B2(n2824), .ZN(
        dp_cluster_3_mult_512_C415_n253) );
  INVD1 U1694 ( .I(dp_cluster_3_mult_513_C415_n86), .ZN(n1260) );
  OAI22D1 U1695 ( .A1(n2685), .A2(n993), .B1(n2809), .B2(n2684), .ZN(
        dp_cluster_3_mult_513_C415_n267) );
  OAI22D1 U1696 ( .A1(n2673), .A2(n2805), .B1(n2806), .B2(n2672), .ZN(
        dp_cluster_3_mult_513_C415_n253) );
  INVD1 U1697 ( .I(dp_cluster_2_mult_486_C409_n86), .ZN(n1258) );
  OAI22D1 U1698 ( .A1(n2359), .A2(n981), .B1(n2483), .B2(n2358), .ZN(
        dp_cluster_2_mult_486_C409_n267) );
  OAI22D1 U1699 ( .A1(n2347), .A2(n2479), .B1(n2480), .B2(n2346), .ZN(
        dp_cluster_2_mult_486_C409_n253) );
  INVD1 U1700 ( .I(dp_cluster_2_mult_485_C409_n86), .ZN(n1117) );
  OAI22D1 U1701 ( .A1(n2511), .A2(n987), .B1(n2635), .B2(n2510), .ZN(
        dp_cluster_2_mult_485_C409_n267) );
  OAI22D1 U1702 ( .A1(n2499), .A2(n2631), .B1(n2632), .B2(n2498), .ZN(
        dp_cluster_2_mult_485_C409_n253) );
  AN2XD1 U1703 ( .A1(n934), .A2(n1148), .Z(n923) );
  AN2XD1 U1704 ( .A1(n923), .A2(n1147), .Z(n924) );
  AN2XD1 U1705 ( .A1(n924), .A2(n1146), .Z(n925) );
  AN2XD1 U1706 ( .A1(n925), .A2(n1145), .Z(n926) );
  AN2XD1 U1707 ( .A1(n926), .A2(n1144), .Z(n927) );
  AN2XD1 U1708 ( .A1(n927), .A2(n1143), .Z(n928) );
  AN2XD1 U1709 ( .A1(n928), .A2(n1142), .Z(n929) );
  AN2XD1 U1710 ( .A1(n929), .A2(n1141), .Z(n930) );
  AN2XD1 U1711 ( .A1(n930), .A2(n1140), .Z(n931) );
  AN2XD1 U1712 ( .A1(n931), .A2(n1139), .Z(n932) );
  AN2XD1 U1713 ( .A1(n932), .A2(n1138), .Z(n933) );
  AN2XD1 U1714 ( .A1(n935), .A2(n1149), .Z(n934) );
  AN2XD1 U1715 ( .A1(n1151), .A2(n1150), .Z(n935) );
  CKXOR2D1 U1716 ( .A1(n1081), .A2(s1_7_i[7]), .Z(n2092) );
  CKXOR2D1 U1717 ( .A1(n1059), .A2(s1_5_i[7]), .Z(n2743) );
  CKXOR2D1 U1718 ( .A1(n1037), .A2(s1_7_r[7]), .Z(n2244) );
  CKXOR2D1 U1719 ( .A1(n1015), .A2(s1_5_r[7]), .Z(n2895) );
  XNR2D1 U1720 ( .A1(n1107), .A2(s1_7_r[3]), .ZN(n1954) );
  XNR2D1 U1721 ( .A1(n1110), .A2(s1_5_r[3]), .ZN(n2605) );
  XNR2D1 U1722 ( .A1(n1101), .A2(s1_7_i[3]), .ZN(n1802) );
  XNR2D1 U1723 ( .A1(n1104), .A2(s1_5_i[3]), .ZN(n2453) );
  XNR2D1 U1724 ( .A1(n1102), .A2(s1_7_i[3]), .ZN(n2128) );
  XNR2D1 U1725 ( .A1(n1105), .A2(s1_5_i[3]), .ZN(n2779) );
  XNR2D1 U1726 ( .A1(n1108), .A2(s1_7_r[3]), .ZN(n2280) );
  XNR2D1 U1727 ( .A1(n1111), .A2(s1_5_r[3]), .ZN(n2931) );
  CKXOR2D1 U1728 ( .A1(n1039), .A2(s1_7_r[5]), .Z(n1936) );
  CKXOR2D1 U1729 ( .A1(n1017), .A2(s1_5_r[5]), .Z(n2587) );
  CKXOR2D1 U1730 ( .A1(n1084), .A2(s1_7_i[5]), .Z(n2110) );
  CKXOR2D1 U1731 ( .A1(n1062), .A2(s1_5_i[5]), .Z(n2761) );
  CKXOR2D1 U1732 ( .A1(n1040), .A2(s1_7_r[5]), .Z(n2262) );
  CKXOR2D1 U1733 ( .A1(n1018), .A2(s1_5_r[5]), .Z(n2913) );
  CKXOR2D1 U1734 ( .A1(n1033), .A2(s1_7_r[9]), .Z(n2304) );
  CKXOR2D1 U1735 ( .A1(n1077), .A2(s1_7_i[9]), .Z(n2152) );
  CKXOR2D1 U1736 ( .A1(n1083), .A2(s1_7_i[5]), .Z(n1784) );
  CKXOR2D1 U1737 ( .A1(n1078), .A2(s1_7_i[9]), .Z(n1826) );
  CKXOR2D1 U1738 ( .A1(n1034), .A2(s1_7_r[9]), .Z(n1978) );
  CKXOR2D1 U1739 ( .A1(n1011), .A2(s1_5_r[9]), .Z(n2955) );
  CKXOR2D1 U1740 ( .A1(n1055), .A2(s1_5_i[9]), .Z(n2803) );
  CKXOR2D1 U1741 ( .A1(n1061), .A2(s1_5_i[5]), .Z(n2435) );
  CKXOR2D1 U1742 ( .A1(n1056), .A2(s1_5_i[9]), .Z(n2477) );
  CKXOR2D1 U1743 ( .A1(n1012), .A2(s1_5_r[9]), .Z(n2629) );
  CKXOR2D1 U1744 ( .A1(n1031), .A2(s1_7_r[11]), .Z(n2300) );
  CKXOR2D1 U1745 ( .A1(n1075), .A2(s1_7_i[11]), .Z(n2148) );
  CKXOR2D1 U1746 ( .A1(n1074), .A2(s1_7_i[11]), .Z(n1822) );
  CKXOR2D1 U1747 ( .A1(n1030), .A2(s1_7_r[11]), .Z(n1974) );
  CKXOR2D1 U1748 ( .A1(n1009), .A2(s1_5_r[11]), .Z(n2951) );
  CKXOR2D1 U1749 ( .A1(n1053), .A2(s1_5_i[11]), .Z(n2799) );
  CKXOR2D1 U1750 ( .A1(n1052), .A2(s1_5_i[11]), .Z(n2473) );
  CKXOR2D1 U1751 ( .A1(n1008), .A2(s1_5_r[11]), .Z(n2625) );
  CKXOR2D1 U1752 ( .A1(n1038), .A2(s1_7_r[7]), .Z(n1918) );
  CKXOR2D1 U1753 ( .A1(n1016), .A2(s1_5_r[7]), .Z(n2569) );
  CKXOR2D1 U1754 ( .A1(n1082), .A2(s1_7_i[7]), .Z(n1766) );
  CKXOR2D1 U1755 ( .A1(n1060), .A2(s1_5_i[7]), .Z(n2417) );
  CKXOR2D1 U1756 ( .A1(n1025), .A2(s1_7_r[15]), .Z(n2307) );
  CKXOR2D1 U1757 ( .A1(n1069), .A2(s1_7_i[15]), .Z(n2155) );
  CKXOR2D1 U1758 ( .A1(n1003), .A2(s1_5_r[15]), .Z(n2958) );
  CKXOR2D1 U1759 ( .A1(n1047), .A2(s1_5_i[15]), .Z(n2806) );
  XNR2D1 U1760 ( .A1(s1_7_r[12]), .A2(s1_7_r[13]), .ZN(n2310) );
  XNR2D1 U1761 ( .A1(s1_5_r[12]), .A2(s1_5_r[13]), .ZN(n2961) );
  XNR2D1 U1762 ( .A1(s1_7_i[12]), .A2(s1_7_i[13]), .ZN(n1832) );
  XNR2D1 U1763 ( .A1(s1_5_i[12]), .A2(s1_5_i[13]), .ZN(n2483) );
  XNR2D1 U1764 ( .A1(s1_7_i[12]), .A2(s1_7_i[13]), .ZN(n2158) );
  XNR2D1 U1765 ( .A1(s1_7_r[12]), .A2(s1_7_r[13]), .ZN(n1984) );
  XNR2D1 U1766 ( .A1(s1_5_i[12]), .A2(s1_5_i[13]), .ZN(n2809) );
  XNR2D1 U1767 ( .A1(s1_5_r[12]), .A2(s1_5_r[13]), .ZN(n2635) );
  CKXOR2D1 U1768 ( .A1(n1026), .A2(s1_7_r[15]), .Z(n1981) );
  CKXOR2D1 U1769 ( .A1(n1004), .A2(s1_5_r[15]), .Z(n2632) );
  CKXOR2D1 U1770 ( .A1(n1070), .A2(s1_7_i[15]), .Z(n1829) );
  CKXOR2D1 U1771 ( .A1(n1048), .A2(s1_5_i[15]), .Z(n2480) );
  NR2D1 U1772 ( .A1(dp_cluster_0_N61), .A2(n1997), .ZN(n1996) );
  OAI22D1 U1773 ( .A1(n1995), .A2(n1171), .B1(dp_cluster_0_N88), .B2(n1994), 
        .ZN(n1997) );
  NR2D1 U1774 ( .A1(dp_cluster_2_N5), .A2(n2648), .ZN(n2647) );
  OAI22D1 U1775 ( .A1(n2646), .A2(n1132), .B1(dp_cluster_2_N32), .B2(n2645), 
        .ZN(n2648) );
  FA1D0 U1776 ( .A(dp_cluster_1_mult_512_C418_n364), .B(
        dp_cluster_1_mult_512_C418_n321), .CI(dp_cluster_1_mult_512_C418_n292), 
        .CO(dp_cluster_1_mult_512_C418_n189), .S(
        dp_cluster_1_mult_512_C418_n190) );
  OAI22D1 U1777 ( .A1(n2284), .A2(n2296), .B1(n2283), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n364) );
  OAI22D1 U1778 ( .A1(n2236), .A2(n974), .B1(n2244), .B2(n2235), .ZN(
        dp_cluster_1_mult_512_C418_n321) );
  OAI22D1 U1779 ( .A1(n2210), .A2(n971), .B1(n2300), .B2(n2209), .ZN(
        dp_cluster_1_mult_512_C418_n292) );
  FA1D0 U1780 ( .A(dp_cluster_1_mult_513_C418_n364), .B(
        dp_cluster_1_mult_513_C418_n321), .CI(dp_cluster_1_mult_513_C418_n292), 
        .CO(dp_cluster_1_mult_513_C418_n189), .S(
        dp_cluster_1_mult_513_C418_n190) );
  OAI22D1 U1781 ( .A1(n2132), .A2(n2144), .B1(n2131), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n364) );
  OAI22D1 U1782 ( .A1(n2084), .A2(n968), .B1(n2092), .B2(n2083), .ZN(
        dp_cluster_1_mult_513_C418_n321) );
  OAI22D1 U1783 ( .A1(n2058), .A2(n965), .B1(n2148), .B2(n2057), .ZN(
        dp_cluster_1_mult_513_C418_n292) );
  FA1D0 U1784 ( .A(dp_cluster_0_mult_486_C412_n364), .B(
        dp_cluster_0_mult_486_C412_n321), .CI(dp_cluster_0_mult_486_C412_n292), 
        .CO(dp_cluster_0_mult_486_C412_n189), .S(
        dp_cluster_0_mult_486_C412_n190) );
  OAI22D1 U1785 ( .A1(n1806), .A2(n1818), .B1(n1805), .B2(n1088), .ZN(
        dp_cluster_0_mult_486_C412_n364) );
  OAI22D1 U1786 ( .A1(n1758), .A2(n956), .B1(n1766), .B2(n1757), .ZN(
        dp_cluster_0_mult_486_C412_n321) );
  OAI22D1 U1787 ( .A1(n1732), .A2(n953), .B1(n1822), .B2(n1731), .ZN(
        dp_cluster_0_mult_486_C412_n292) );
  FA1D0 U1788 ( .A(dp_cluster_0_mult_485_C412_n364), .B(
        dp_cluster_0_mult_485_C412_n321), .CI(dp_cluster_0_mult_485_C412_n292), 
        .CO(dp_cluster_0_mult_485_C412_n189), .S(
        dp_cluster_0_mult_485_C412_n190) );
  OAI22D1 U1789 ( .A1(n1958), .A2(n1970), .B1(n1957), .B2(n1044), .ZN(
        dp_cluster_0_mult_485_C412_n364) );
  OAI22D1 U1790 ( .A1(n1910), .A2(n962), .B1(n1918), .B2(n1909), .ZN(
        dp_cluster_0_mult_485_C412_n321) );
  OAI22D1 U1791 ( .A1(n1884), .A2(n959), .B1(n1974), .B2(n1883), .ZN(
        dp_cluster_0_mult_485_C412_n292) );
  FA1D0 U1792 ( .A(dp_cluster_3_mult_512_C415_n364), .B(
        dp_cluster_3_mult_512_C415_n321), .CI(dp_cluster_3_mult_512_C415_n292), 
        .CO(dp_cluster_3_mult_512_C415_n189), .S(
        dp_cluster_3_mult_512_C415_n190) );
  OAI22D1 U1793 ( .A1(n2935), .A2(n2947), .B1(n2934), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n364) );
  OAI22D1 U1794 ( .A1(n2887), .A2(n998), .B1(n2895), .B2(n2886), .ZN(
        dp_cluster_3_mult_512_C415_n321) );
  OAI22D1 U1795 ( .A1(n2861), .A2(n995), .B1(n2951), .B2(n2860), .ZN(
        dp_cluster_3_mult_512_C415_n292) );
  FA1D0 U1796 ( .A(dp_cluster_3_mult_513_C415_n364), .B(
        dp_cluster_3_mult_513_C415_n321), .CI(dp_cluster_3_mult_513_C415_n292), 
        .CO(dp_cluster_3_mult_513_C415_n189), .S(
        dp_cluster_3_mult_513_C415_n190) );
  OAI22D1 U1797 ( .A1(n2783), .A2(n2795), .B1(n2782), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n364) );
  OAI22D1 U1798 ( .A1(n2735), .A2(n992), .B1(n2743), .B2(n2734), .ZN(
        dp_cluster_3_mult_513_C415_n321) );
  OAI22D1 U1799 ( .A1(n2709), .A2(n989), .B1(n2799), .B2(n2708), .ZN(
        dp_cluster_3_mult_513_C415_n292) );
  FA1D0 U1800 ( .A(dp_cluster_2_mult_486_C409_n364), .B(
        dp_cluster_2_mult_486_C409_n321), .CI(dp_cluster_2_mult_486_C409_n292), 
        .CO(dp_cluster_2_mult_486_C409_n189), .S(
        dp_cluster_2_mult_486_C409_n190) );
  OAI22D1 U1801 ( .A1(n2457), .A2(n2469), .B1(n2456), .B2(n1066), .ZN(
        dp_cluster_2_mult_486_C409_n364) );
  OAI22D1 U1802 ( .A1(n2409), .A2(n980), .B1(n2417), .B2(n2408), .ZN(
        dp_cluster_2_mult_486_C409_n321) );
  OAI22D1 U1803 ( .A1(n2383), .A2(n977), .B1(n2473), .B2(n2382), .ZN(
        dp_cluster_2_mult_486_C409_n292) );
  FA1D0 U1804 ( .A(dp_cluster_2_mult_485_C409_n364), .B(
        dp_cluster_2_mult_485_C409_n321), .CI(dp_cluster_2_mult_485_C409_n292), 
        .CO(dp_cluster_2_mult_485_C409_n189), .S(
        dp_cluster_2_mult_485_C409_n190) );
  OAI22D1 U1805 ( .A1(n2609), .A2(n2621), .B1(n2608), .B2(n1022), .ZN(
        dp_cluster_2_mult_485_C409_n364) );
  OAI22D1 U1806 ( .A1(n2561), .A2(n986), .B1(n2569), .B2(n2560), .ZN(
        dp_cluster_2_mult_485_C409_n321) );
  OAI22D1 U1807 ( .A1(n2535), .A2(n983), .B1(n2625), .B2(n2534), .ZN(
        dp_cluster_2_mult_485_C409_n292) );
  INVD1 U1808 ( .I(s1_7_r[10]), .ZN(n1163) );
  INVD1 U1809 ( .I(s1_5_r[10]), .ZN(n1124) );
  INVD1 U1810 ( .I(s1_7_i[14]), .ZN(n1288) );
  INVD1 U1811 ( .I(s1_7_r[14]), .ZN(n1153) );
  INVD1 U1812 ( .I(s1_5_i[14]), .ZN(n1255) );
  INVD1 U1813 ( .I(s1_5_r[14]), .ZN(n1114) );
  INVD1 U1814 ( .I(s1_7_r[4]), .ZN(n1173) );
  INVD1 U1815 ( .I(s1_5_r[4]), .ZN(n1134) );
  INVD1 U1816 ( .I(s1_7_r[6]), .ZN(n1169) );
  INVD1 U1817 ( .I(s1_5_r[6]), .ZN(n1130) );
  INVD1 U1818 ( .I(s1_7_i[4]), .ZN(n1304) );
  INVD1 U1819 ( .I(s1_5_i[4]), .ZN(n1271) );
  INVD1 U1820 ( .I(s1_7_i[6]), .ZN(n1301) );
  INVD1 U1821 ( .I(s1_5_i[6]), .ZN(n1268) );
  INVD1 U1822 ( .I(s1_7_r[8]), .ZN(n1165) );
  INVD1 U1823 ( .I(s1_7_i[8]), .ZN(n1298) );
  INVD1 U1824 ( .I(s1_5_r[8]), .ZN(n1126) );
  INVD1 U1825 ( .I(s1_5_i[8]), .ZN(n1265) );
  INVD1 U1826 ( .I(s1_7_i[10]), .ZN(n1297) );
  INVD1 U1827 ( .I(s1_5_i[10]), .ZN(n1264) );
  INVD1 U1828 ( .I(s1_7_r[1]), .ZN(n1175) );
  INVD1 U1829 ( .I(s1_5_r[1]), .ZN(n1136) );
  INVD1 U1830 ( .I(s1_7_i[1]), .ZN(n1305) );
  INVD1 U1831 ( .I(s1_5_i[1]), .ZN(n1272) );
  OAI22D1 U1832 ( .A1(n2193), .A2(n975), .B1(n2310), .B2(n2192), .ZN(
        dp_cluster_1_mult_512_C418_n274) );
  OAI22D1 U1833 ( .A1(n2181), .A2(n2306), .B1(n2307), .B2(n2180), .ZN(
        dp_cluster_1_mult_512_C418_n260) );
  OAI22D1 U1834 ( .A1(n2041), .A2(n969), .B1(n2158), .B2(n2040), .ZN(
        dp_cluster_1_mult_513_C418_n274) );
  OAI22D1 U1835 ( .A1(n2029), .A2(n2154), .B1(n2155), .B2(n2028), .ZN(
        dp_cluster_1_mult_513_C418_n260) );
  OAI22D1 U1836 ( .A1(n2844), .A2(n999), .B1(n2961), .B2(n2843), .ZN(
        dp_cluster_3_mult_512_C415_n274) );
  OAI22D1 U1837 ( .A1(n2832), .A2(n2957), .B1(n2958), .B2(n2831), .ZN(
        dp_cluster_3_mult_512_C415_n260) );
  OAI22D1 U1838 ( .A1(n2692), .A2(n993), .B1(n2809), .B2(n2691), .ZN(
        dp_cluster_3_mult_513_C415_n274) );
  OAI22D1 U1839 ( .A1(n2680), .A2(n2805), .B1(n2806), .B2(n2679), .ZN(
        dp_cluster_3_mult_513_C415_n260) );
  ND2D1 U1840 ( .A1(n2307), .A2(n2171), .ZN(n2306) );
  ND2D1 U1841 ( .A1(n2155), .A2(n2019), .ZN(n2154) );
  ND2D1 U1842 ( .A1(n2958), .A2(n2822), .ZN(n2957) );
  ND2D1 U1843 ( .A1(n2806), .A2(n2670), .ZN(n2805) );
  ND2D1 U1844 ( .A1(n1981), .A2(n1845), .ZN(n1980) );
  ND2D1 U1845 ( .A1(n2632), .A2(n2496), .ZN(n2631) );
  ND2D1 U1846 ( .A1(n1829), .A2(n1693), .ZN(n1828) );
  ND2D1 U1847 ( .A1(n2480), .A2(n2344), .ZN(n2479) );
  INVD1 U1848 ( .I(s1_7_i[12]), .ZN(n1294) );
  INVD1 U1849 ( .I(s1_7_r[12]), .ZN(n1159) );
  INVD1 U1850 ( .I(s1_5_i[12]), .ZN(n1261) );
  INVD1 U1851 ( .I(s1_5_r[12]), .ZN(n1120) );
  CKBD1 U1852 ( .I(n1934), .Z(n960) );
  ND2D1 U1853 ( .A1(n1936), .A2(n1839), .ZN(n1934) );
  CKBD1 U1854 ( .I(n2585), .Z(n984) );
  ND2D1 U1855 ( .A1(n2587), .A2(n2490), .ZN(n2585) );
  CKBD1 U1856 ( .I(n2108), .Z(n966) );
  ND2D1 U1857 ( .A1(n2110), .A2(n2013), .ZN(n2108) );
  CKBD1 U1858 ( .I(n2126), .Z(n967) );
  ND2D1 U1859 ( .A1(n2128), .A2(n2014), .ZN(n2126) );
  CKBD1 U1860 ( .I(n2759), .Z(n990) );
  ND2D1 U1861 ( .A1(n2761), .A2(n2664), .ZN(n2759) );
  CKBD1 U1862 ( .I(n2777), .Z(n991) );
  ND2D1 U1863 ( .A1(n2779), .A2(n2665), .ZN(n2777) );
  CKBD1 U1864 ( .I(n2090), .Z(n968) );
  ND2D1 U1865 ( .A1(n2092), .A2(n2015), .ZN(n2090) );
  CKBD1 U1866 ( .I(n1916), .Z(n962) );
  ND2D1 U1867 ( .A1(n1918), .A2(n1841), .ZN(n1916) );
  CKBD1 U1868 ( .I(n2741), .Z(n992) );
  ND2D1 U1869 ( .A1(n2743), .A2(n2666), .ZN(n2741) );
  CKBD1 U1870 ( .I(n2567), .Z(n986) );
  ND2D1 U1871 ( .A1(n2569), .A2(n2492), .ZN(n2567) );
  CKBD1 U1872 ( .I(n2242), .Z(n974) );
  ND2D1 U1873 ( .A1(n2244), .A2(n2167), .ZN(n2242) );
  CKBD1 U1874 ( .I(n2260), .Z(n972) );
  ND2D1 U1875 ( .A1(n2262), .A2(n2165), .ZN(n2260) );
  CKBD1 U1876 ( .I(n2278), .Z(n973) );
  ND2D1 U1877 ( .A1(n2280), .A2(n2166), .ZN(n2278) );
  CKBD1 U1878 ( .I(n2893), .Z(n998) );
  ND2D1 U1879 ( .A1(n2895), .A2(n2818), .ZN(n2893) );
  CKBD1 U1880 ( .I(n2911), .Z(n996) );
  ND2D1 U1881 ( .A1(n2913), .A2(n2816), .ZN(n2911) );
  CKBD1 U1882 ( .I(n2929), .Z(n997) );
  ND2D1 U1883 ( .A1(n2931), .A2(n2817), .ZN(n2929) );
  CKBD1 U1884 ( .I(n2301), .Z(n976) );
  ND2D1 U1885 ( .A1(n2304), .A2(n2172), .ZN(n2301) );
  CKBD1 U1886 ( .I(n2149), .Z(n970) );
  ND2D1 U1887 ( .A1(n2152), .A2(n2020), .ZN(n2149) );
  CKBD1 U1888 ( .I(n1764), .Z(n956) );
  ND2D1 U1889 ( .A1(n1766), .A2(n1689), .ZN(n1764) );
  CKBD1 U1890 ( .I(n1782), .Z(n954) );
  ND2D1 U1891 ( .A1(n1784), .A2(n1687), .ZN(n1782) );
  CKBD1 U1892 ( .I(n1823), .Z(n958) );
  ND2D1 U1893 ( .A1(n1826), .A2(n1694), .ZN(n1823) );
  CKBD1 U1894 ( .I(n1975), .Z(n964) );
  ND2D1 U1895 ( .A1(n1978), .A2(n1846), .ZN(n1975) );
  CKBD1 U1896 ( .I(n2952), .Z(n1000) );
  ND2D1 U1897 ( .A1(n2955), .A2(n2823), .ZN(n2952) );
  CKBD1 U1898 ( .I(n2800), .Z(n994) );
  ND2D1 U1899 ( .A1(n2803), .A2(n2671), .ZN(n2800) );
  CKBD1 U1900 ( .I(n2415), .Z(n980) );
  ND2D1 U1901 ( .A1(n2417), .A2(n2340), .ZN(n2415) );
  CKBD1 U1902 ( .I(n2433), .Z(n978) );
  ND2D1 U1903 ( .A1(n2435), .A2(n2338), .ZN(n2433) );
  CKBD1 U1904 ( .I(n2474), .Z(n982) );
  ND2D1 U1905 ( .A1(n2477), .A2(n2345), .ZN(n2474) );
  CKBD1 U1906 ( .I(n2626), .Z(n988) );
  ND2D1 U1907 ( .A1(n2629), .A2(n2497), .ZN(n2626) );
  CKBD1 U1908 ( .I(n2311), .Z(n975) );
  ND2D1 U1909 ( .A1(n2310), .A2(n2168), .ZN(n2311) );
  CKBD1 U1910 ( .I(n2297), .Z(n971) );
  ND2D1 U1911 ( .A1(n2300), .A2(n2164), .ZN(n2297) );
  CKBD1 U1912 ( .I(n2145), .Z(n965) );
  ND2D1 U1913 ( .A1(n2148), .A2(n2012), .ZN(n2145) );
  CKBD1 U1914 ( .I(n1819), .Z(n953) );
  ND2D1 U1915 ( .A1(n1822), .A2(n1686), .ZN(n1819) );
  CKBD1 U1916 ( .I(n1971), .Z(n959) );
  ND2D1 U1917 ( .A1(n1974), .A2(n1838), .ZN(n1971) );
  CKBD1 U1918 ( .I(n2962), .Z(n999) );
  ND2D1 U1919 ( .A1(n2961), .A2(n2819), .ZN(n2962) );
  CKBD1 U1920 ( .I(n2948), .Z(n995) );
  ND2D1 U1921 ( .A1(n2951), .A2(n2815), .ZN(n2948) );
  CKBD1 U1922 ( .I(n2796), .Z(n989) );
  ND2D1 U1923 ( .A1(n2799), .A2(n2663), .ZN(n2796) );
  CKBD1 U1924 ( .I(n2470), .Z(n977) );
  ND2D1 U1925 ( .A1(n2473), .A2(n2337), .ZN(n2470) );
  CKBD1 U1926 ( .I(n2622), .Z(n983) );
  ND2D1 U1927 ( .A1(n2625), .A2(n2489), .ZN(n2622) );
  CKBD1 U1928 ( .I(n1833), .Z(n957) );
  ND2D1 U1929 ( .A1(n1832), .A2(n1690), .ZN(n1833) );
  CKBD1 U1930 ( .I(n2484), .Z(n981) );
  ND2D1 U1931 ( .A1(n2483), .A2(n2341), .ZN(n2484) );
  CKBD1 U1932 ( .I(n2159), .Z(n969) );
  ND2D1 U1933 ( .A1(n2158), .A2(n2016), .ZN(n2159) );
  CKBD1 U1934 ( .I(n1985), .Z(n963) );
  ND2D1 U1935 ( .A1(n1984), .A2(n1842), .ZN(n1985) );
  CKBD1 U1936 ( .I(n2810), .Z(n993) );
  ND2D1 U1937 ( .A1(n2809), .A2(n2667), .ZN(n2810) );
  CKBD1 U1938 ( .I(n2636), .Z(n987) );
  ND2D1 U1939 ( .A1(n2635), .A2(n2493), .ZN(n2636) );
  INVD1 U1940 ( .I(s1_7_i[16]), .ZN(n1285) );
  INVD1 U1941 ( .I(s1_7_r[16]), .ZN(n1152) );
  INVD1 U1942 ( .I(s1_5_i[16]), .ZN(n1252) );
  INVD1 U1943 ( .I(s1_5_r[16]), .ZN(n1113) );
  OAI22D1 U1944 ( .A1(n1965), .A2(n1970), .B1(n1964), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n371) );
  OAI22D1 U1945 ( .A1(n1949), .A2(n961), .B1(n1954), .B2(n1948), .ZN(
        dp_cluster_0_mult_485_C412_n356) );
  NR2D1 U1946 ( .A1(n1918), .A2(n1093), .ZN(dp_cluster_0_mult_485_C412_n328)
         );
  OAI22D1 U1947 ( .A1(n2616), .A2(n2621), .B1(n2615), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n371) );
  OAI22D1 U1948 ( .A1(n2600), .A2(n985), .B1(n2605), .B2(n2599), .ZN(
        dp_cluster_2_mult_485_C409_n356) );
  NR2D1 U1949 ( .A1(n2569), .A2(n1090), .ZN(dp_cluster_2_mult_485_C409_n328)
         );
  OAI22D1 U1950 ( .A1(n2137), .A2(n2144), .B1(n2136), .B2(n1087), .ZN(
        dp_cluster_1_mult_513_C418_n369) );
  OAI22D1 U1951 ( .A1(n2121), .A2(n967), .B1(n2128), .B2(n2120), .ZN(
        dp_cluster_1_mult_513_C418_n354) );
  OAI22D1 U1952 ( .A1(n1963), .A2(n1970), .B1(n1962), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n369) );
  OAI22D1 U1953 ( .A1(n1947), .A2(n961), .B1(n1954), .B2(n1946), .ZN(
        dp_cluster_0_mult_485_C412_n354) );
  OAI22D1 U1954 ( .A1(n2788), .A2(n2795), .B1(n2787), .B2(n1065), .ZN(
        dp_cluster_3_mult_513_C415_n369) );
  OAI22D1 U1955 ( .A1(n2772), .A2(n991), .B1(n2779), .B2(n2771), .ZN(
        dp_cluster_3_mult_513_C415_n354) );
  OAI22D1 U1956 ( .A1(n2614), .A2(n2621), .B1(n2613), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n369) );
  OAI22D1 U1957 ( .A1(n2598), .A2(n985), .B1(n2605), .B2(n2597), .ZN(
        dp_cluster_2_mult_485_C409_n354) );
  OAI22D1 U1958 ( .A1(n2136), .A2(n2144), .B1(n2135), .B2(n1087), .ZN(
        dp_cluster_1_mult_513_C418_n368) );
  OAI22D1 U1959 ( .A1(n1962), .A2(n1970), .B1(n1961), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n368) );
  OAI22D1 U1960 ( .A1(n2787), .A2(n2795), .B1(n2786), .B2(n1065), .ZN(
        dp_cluster_3_mult_513_C415_n368) );
  OAI22D1 U1961 ( .A1(n2613), .A2(n2621), .B1(n2612), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n368) );
  OAI22D1 U1962 ( .A1(n2135), .A2(n2144), .B1(n2134), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n367) );
  OAI22D1 U1963 ( .A1(n2119), .A2(n967), .B1(n2128), .B2(n2118), .ZN(
        dp_cluster_1_mult_513_C418_n352) );
  OAI22D1 U1964 ( .A1(n1961), .A2(n1970), .B1(n1960), .B2(n1044), .ZN(
        dp_cluster_0_mult_485_C412_n367) );
  OAI22D1 U1965 ( .A1(n1945), .A2(n961), .B1(n1954), .B2(n1944), .ZN(
        dp_cluster_0_mult_485_C412_n352) );
  OAI22D1 U1966 ( .A1(n2786), .A2(n2795), .B1(n2785), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n367) );
  OAI22D1 U1967 ( .A1(n2770), .A2(n991), .B1(n2779), .B2(n2769), .ZN(
        dp_cluster_3_mult_513_C415_n352) );
  OAI22D1 U1968 ( .A1(n2612), .A2(n2621), .B1(n2611), .B2(n1022), .ZN(
        dp_cluster_2_mult_485_C409_n367) );
  OAI22D1 U1969 ( .A1(n2596), .A2(n985), .B1(n2605), .B2(n2595), .ZN(
        dp_cluster_2_mult_485_C409_n352) );
  OAI22D1 U1970 ( .A1(n2238), .A2(n974), .B1(n2244), .B2(n2237), .ZN(
        dp_cluster_1_mult_512_C418_n323) );
  OAI22D1 U1971 ( .A1(n2086), .A2(n968), .B1(n2092), .B2(n2085), .ZN(
        dp_cluster_1_mult_513_C418_n323) );
  OAI22D1 U1972 ( .A1(n1912), .A2(n962), .B1(n1918), .B2(n1911), .ZN(
        dp_cluster_0_mult_485_C412_n323) );
  OAI22D1 U1973 ( .A1(n2889), .A2(n998), .B1(n2895), .B2(n2888), .ZN(
        dp_cluster_3_mult_512_C415_n323) );
  OAI22D1 U1974 ( .A1(n2737), .A2(n992), .B1(n2743), .B2(n2736), .ZN(
        dp_cluster_3_mult_513_C415_n323) );
  OAI22D1 U1975 ( .A1(n2563), .A2(n986), .B1(n2569), .B2(n2562), .ZN(
        dp_cluster_2_mult_485_C409_n323) );
  OAI22D1 U1976 ( .A1(n2221), .A2(n976), .B1(n2304), .B2(n2220), .ZN(
        dp_cluster_1_mult_512_C418_n305) );
  OAI22D1 U1977 ( .A1(n2209), .A2(n971), .B1(n2300), .B2(n2208), .ZN(
        dp_cluster_1_mult_512_C418_n291) );
  NR2D1 U1978 ( .A1(n2307), .A2(n1099), .ZN(dp_cluster_1_mult_512_C418_n264)
         );
  OAI22D1 U1979 ( .A1(n2069), .A2(n970), .B1(n2152), .B2(n2068), .ZN(
        dp_cluster_1_mult_513_C418_n305) );
  OAI22D1 U1980 ( .A1(n2057), .A2(n965), .B1(n2148), .B2(n2056), .ZN(
        dp_cluster_1_mult_513_C418_n291) );
  NR2D1 U1981 ( .A1(n2155), .A2(n1093), .ZN(dp_cluster_1_mult_513_C418_n264)
         );
  OAI22D1 U1982 ( .A1(n1743), .A2(n958), .B1(n1826), .B2(n1742), .ZN(
        dp_cluster_0_mult_486_C412_n305) );
  OAI22D1 U1983 ( .A1(n1731), .A2(n953), .B1(n1822), .B2(n1730), .ZN(
        dp_cluster_0_mult_486_C412_n291) );
  NR2D1 U1984 ( .A1(n1829), .A2(n1100), .ZN(dp_cluster_0_mult_486_C412_n264)
         );
  OAI22D1 U1985 ( .A1(n1895), .A2(n964), .B1(n1978), .B2(n1894), .ZN(
        dp_cluster_0_mult_485_C412_n305) );
  OAI22D1 U1986 ( .A1(n1883), .A2(n959), .B1(n1974), .B2(n1882), .ZN(
        dp_cluster_0_mult_485_C412_n291) );
  NR2D1 U1987 ( .A1(n1981), .A2(n1094), .ZN(dp_cluster_0_mult_485_C412_n264)
         );
  OAI22D1 U1988 ( .A1(n2872), .A2(n1000), .B1(n2955), .B2(n2871), .ZN(
        dp_cluster_3_mult_512_C415_n305) );
  OAI22D1 U1989 ( .A1(n2860), .A2(n995), .B1(n2951), .B2(n2859), .ZN(
        dp_cluster_3_mult_512_C415_n291) );
  NR2D1 U1990 ( .A1(n2958), .A2(n1096), .ZN(dp_cluster_3_mult_512_C415_n264)
         );
  OAI22D1 U1991 ( .A1(n2720), .A2(n994), .B1(n2803), .B2(n2719), .ZN(
        dp_cluster_3_mult_513_C415_n305) );
  OAI22D1 U1992 ( .A1(n2708), .A2(n989), .B1(n2799), .B2(n2707), .ZN(
        dp_cluster_3_mult_513_C415_n291) );
  NR2D1 U1993 ( .A1(n2806), .A2(n1090), .ZN(dp_cluster_3_mult_513_C415_n264)
         );
  OAI22D1 U1994 ( .A1(n2394), .A2(n982), .B1(n2477), .B2(n2393), .ZN(
        dp_cluster_2_mult_486_C409_n305) );
  OAI22D1 U1995 ( .A1(n2382), .A2(n977), .B1(n2473), .B2(n2381), .ZN(
        dp_cluster_2_mult_486_C409_n291) );
  NR2D1 U1996 ( .A1(n2480), .A2(n1097), .ZN(dp_cluster_2_mult_486_C409_n264)
         );
  OAI22D1 U1997 ( .A1(n2546), .A2(n988), .B1(n2629), .B2(n2545), .ZN(
        dp_cluster_2_mult_485_C409_n305) );
  OAI22D1 U1998 ( .A1(n2534), .A2(n983), .B1(n2625), .B2(n2533), .ZN(
        dp_cluster_2_mult_485_C409_n291) );
  NR2D1 U1999 ( .A1(n2632), .A2(n1091), .ZN(dp_cluster_2_mult_485_C409_n264)
         );
  OAI22D1 U2000 ( .A1(n2234), .A2(n974), .B1(n2244), .B2(n2233), .ZN(
        dp_cluster_1_mult_512_C418_n319) );
  OAI22D1 U2001 ( .A1(n2208), .A2(n971), .B1(n2300), .B2(n2207), .ZN(
        dp_cluster_1_mult_512_C418_n290) );
  OAI22D1 U2002 ( .A1(n2196), .A2(n975), .B1(n2310), .B2(n2195), .ZN(
        dp_cluster_1_mult_512_C418_n277) );
  OAI22D1 U2003 ( .A1(n2082), .A2(n968), .B1(n2092), .B2(n2081), .ZN(
        dp_cluster_1_mult_513_C418_n319) );
  OAI22D1 U2004 ( .A1(n2056), .A2(n965), .B1(n2148), .B2(n2055), .ZN(
        dp_cluster_1_mult_513_C418_n290) );
  OAI22D1 U2005 ( .A1(n2044), .A2(n969), .B1(n2158), .B2(n2043), .ZN(
        dp_cluster_1_mult_513_C418_n277) );
  OAI22D1 U2006 ( .A1(n1756), .A2(n956), .B1(n1766), .B2(n1755), .ZN(
        dp_cluster_0_mult_486_C412_n319) );
  OAI22D1 U2007 ( .A1(n1730), .A2(n953), .B1(n1822), .B2(n1729), .ZN(
        dp_cluster_0_mult_486_C412_n290) );
  OAI22D1 U2008 ( .A1(n1718), .A2(n957), .B1(n1832), .B2(n1717), .ZN(
        dp_cluster_0_mult_486_C412_n277) );
  OAI22D1 U2009 ( .A1(n1908), .A2(n962), .B1(n1918), .B2(n1907), .ZN(
        dp_cluster_0_mult_485_C412_n319) );
  OAI22D1 U2010 ( .A1(n1882), .A2(n959), .B1(n1974), .B2(n1881), .ZN(
        dp_cluster_0_mult_485_C412_n290) );
  OAI22D1 U2011 ( .A1(n1870), .A2(n963), .B1(n1984), .B2(n1869), .ZN(
        dp_cluster_0_mult_485_C412_n277) );
  OAI22D1 U2012 ( .A1(n2885), .A2(n998), .B1(n2895), .B2(n2884), .ZN(
        dp_cluster_3_mult_512_C415_n319) );
  OAI22D1 U2013 ( .A1(n2859), .A2(n995), .B1(n2951), .B2(n2858), .ZN(
        dp_cluster_3_mult_512_C415_n290) );
  OAI22D1 U2014 ( .A1(n2847), .A2(n999), .B1(n2961), .B2(n2846), .ZN(
        dp_cluster_3_mult_512_C415_n277) );
  OAI22D1 U2015 ( .A1(n2733), .A2(n992), .B1(n2743), .B2(n2732), .ZN(
        dp_cluster_3_mult_513_C415_n319) );
  OAI22D1 U2016 ( .A1(n2707), .A2(n989), .B1(n2799), .B2(n2706), .ZN(
        dp_cluster_3_mult_513_C415_n290) );
  OAI22D1 U2017 ( .A1(n2695), .A2(n993), .B1(n2809), .B2(n2694), .ZN(
        dp_cluster_3_mult_513_C415_n277) );
  OAI22D1 U2018 ( .A1(n2407), .A2(n980), .B1(n2417), .B2(n2406), .ZN(
        dp_cluster_2_mult_486_C409_n319) );
  OAI22D1 U2019 ( .A1(n2381), .A2(n977), .B1(n2473), .B2(n2380), .ZN(
        dp_cluster_2_mult_486_C409_n290) );
  OAI22D1 U2020 ( .A1(n2369), .A2(n981), .B1(n2483), .B2(n2368), .ZN(
        dp_cluster_2_mult_486_C409_n277) );
  OAI22D1 U2021 ( .A1(n2559), .A2(n986), .B1(n2569), .B2(n2558), .ZN(
        dp_cluster_2_mult_485_C409_n319) );
  OAI22D1 U2022 ( .A1(n2533), .A2(n983), .B1(n2625), .B2(n2532), .ZN(
        dp_cluster_2_mult_485_C409_n290) );
  OAI22D1 U2023 ( .A1(n2521), .A2(n987), .B1(n2635), .B2(n2520), .ZN(
        dp_cluster_2_mult_485_C409_n277) );
  OAI22D1 U2024 ( .A1(n1715), .A2(n957), .B1(n1832), .B2(n1714), .ZN(
        dp_cluster_0_mult_486_C412_n274) );
  OAI22D1 U2025 ( .A1(n1703), .A2(n1828), .B1(n1829), .B2(n1702), .ZN(
        dp_cluster_0_mult_486_C412_n260) );
  OAI22D1 U2026 ( .A1(n1867), .A2(n963), .B1(n1984), .B2(n1866), .ZN(
        dp_cluster_0_mult_485_C412_n274) );
  OAI22D1 U2027 ( .A1(n1855), .A2(n1980), .B1(n1981), .B2(n1854), .ZN(
        dp_cluster_0_mult_485_C412_n260) );
  OAI22D1 U2028 ( .A1(n2366), .A2(n981), .B1(n2483), .B2(n2365), .ZN(
        dp_cluster_2_mult_486_C409_n274) );
  OAI22D1 U2029 ( .A1(n2354), .A2(n2479), .B1(n2480), .B2(n2353), .ZN(
        dp_cluster_2_mult_486_C409_n260) );
  OAI22D1 U2030 ( .A1(n2518), .A2(n987), .B1(n2635), .B2(n2517), .ZN(
        dp_cluster_2_mult_485_C409_n274) );
  OAI22D1 U2031 ( .A1(n2506), .A2(n2631), .B1(n2632), .B2(n2505), .ZN(
        dp_cluster_2_mult_485_C409_n260) );
  OAI22D1 U2032 ( .A1(n2139), .A2(n2144), .B1(n2138), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n371) );
  OAI22D1 U2033 ( .A1(n2123), .A2(n967), .B1(n2128), .B2(n2122), .ZN(
        dp_cluster_1_mult_513_C418_n356) );
  NR2D1 U2034 ( .A1(n2092), .A2(n1092), .ZN(dp_cluster_1_mult_513_C418_n328)
         );
  OAI22D1 U2035 ( .A1(n2790), .A2(n2795), .B1(n2789), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n371) );
  OAI22D1 U2036 ( .A1(n2774), .A2(n991), .B1(n2779), .B2(n2773), .ZN(
        dp_cluster_3_mult_513_C415_n356) );
  NR2D1 U2037 ( .A1(n2743), .A2(n1089), .ZN(dp_cluster_3_mult_513_C415_n328)
         );
  OAI22D1 U2038 ( .A1(n2291), .A2(n2296), .B1(n2290), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n371) );
  OAI22D1 U2039 ( .A1(n2275), .A2(n973), .B1(n2280), .B2(n2274), .ZN(
        dp_cluster_1_mult_512_C418_n356) );
  NR2D1 U2040 ( .A1(n2244), .A2(n1098), .ZN(dp_cluster_1_mult_512_C418_n328)
         );
  OAI22D1 U2041 ( .A1(n2942), .A2(n2947), .B1(n2941), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n371) );
  OAI22D1 U2042 ( .A1(n2926), .A2(n997), .B1(n2931), .B2(n2925), .ZN(
        dp_cluster_3_mult_512_C415_n356) );
  NR2D1 U2043 ( .A1(n2895), .A2(n1095), .ZN(dp_cluster_3_mult_512_C415_n328)
         );
  OAI22D1 U2044 ( .A1(n1813), .A2(n1818), .B1(n1812), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n371) );
  OAI22D1 U2045 ( .A1(n1797), .A2(n955), .B1(n1802), .B2(n1796), .ZN(
        dp_cluster_0_mult_486_C412_n356) );
  NR2D1 U2046 ( .A1(n1766), .A2(n1099), .ZN(dp_cluster_0_mult_486_C412_n328)
         );
  OAI22D1 U2047 ( .A1(n2464), .A2(n2469), .B1(n2463), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n371) );
  OAI22D1 U2048 ( .A1(n2448), .A2(n979), .B1(n2453), .B2(n2447), .ZN(
        dp_cluster_2_mult_486_C409_n356) );
  NR2D1 U2049 ( .A1(n2417), .A2(n1096), .ZN(dp_cluster_2_mult_486_C409_n328)
         );
  OAI22D1 U2050 ( .A1(n2289), .A2(n2296), .B1(n2288), .B2(n1043), .ZN(
        dp_cluster_1_mult_512_C418_n369) );
  OAI22D1 U2051 ( .A1(n2273), .A2(n973), .B1(n2280), .B2(n2272), .ZN(
        dp_cluster_1_mult_512_C418_n354) );
  OAI22D1 U2052 ( .A1(n1811), .A2(n1818), .B1(n1810), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n369) );
  OAI22D1 U2053 ( .A1(n1795), .A2(n955), .B1(n1802), .B2(n1794), .ZN(
        dp_cluster_0_mult_486_C412_n354) );
  OAI22D1 U2054 ( .A1(n2940), .A2(n2947), .B1(n2939), .B2(n1021), .ZN(
        dp_cluster_3_mult_512_C415_n369) );
  OAI22D1 U2055 ( .A1(n2924), .A2(n997), .B1(n2931), .B2(n2923), .ZN(
        dp_cluster_3_mult_512_C415_n354) );
  OAI22D1 U2056 ( .A1(n2462), .A2(n2469), .B1(n2461), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n369) );
  OAI22D1 U2057 ( .A1(n2446), .A2(n979), .B1(n2453), .B2(n2445), .ZN(
        dp_cluster_2_mult_486_C409_n354) );
  OAI22D1 U2058 ( .A1(n2288), .A2(n2296), .B1(n2287), .B2(n1043), .ZN(
        dp_cluster_1_mult_512_C418_n368) );
  OAI22D1 U2059 ( .A1(n1810), .A2(n1818), .B1(n1809), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n368) );
  OAI22D1 U2060 ( .A1(n2939), .A2(n2947), .B1(n2938), .B2(n1021), .ZN(
        dp_cluster_3_mult_512_C415_n368) );
  OAI22D1 U2061 ( .A1(n2461), .A2(n2469), .B1(n2460), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n368) );
  OAI22D1 U2062 ( .A1(n2287), .A2(n2296), .B1(n2286), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n367) );
  OAI22D1 U2063 ( .A1(n2271), .A2(n973), .B1(n2280), .B2(n2270), .ZN(
        dp_cluster_1_mult_512_C418_n352) );
  OAI22D1 U2064 ( .A1(n1809), .A2(n1818), .B1(n1808), .B2(n1088), .ZN(
        dp_cluster_0_mult_486_C412_n367) );
  OAI22D1 U2065 ( .A1(n1793), .A2(n955), .B1(n1802), .B2(n1792), .ZN(
        dp_cluster_0_mult_486_C412_n352) );
  OAI22D1 U2066 ( .A1(n2938), .A2(n2947), .B1(n2937), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n367) );
  OAI22D1 U2067 ( .A1(n2922), .A2(n997), .B1(n2931), .B2(n2921), .ZN(
        dp_cluster_3_mult_512_C415_n352) );
  OAI22D1 U2068 ( .A1(n2460), .A2(n2469), .B1(n2459), .B2(n1066), .ZN(
        dp_cluster_2_mult_486_C409_n367) );
  OAI22D1 U2069 ( .A1(n2444), .A2(n979), .B1(n2453), .B2(n2443), .ZN(
        dp_cluster_2_mult_486_C409_n352) );
  OAI22D1 U2070 ( .A1(n1760), .A2(n956), .B1(n1766), .B2(n1759), .ZN(
        dp_cluster_0_mult_486_C412_n323) );
  OAI22D1 U2071 ( .A1(n2411), .A2(n980), .B1(n2417), .B2(n2410), .ZN(
        dp_cluster_2_mult_486_C409_n323) );
  FA1D0 U2072 ( .A(dp_cluster_0_mult_485_C412_n373), .B(
        dp_cluster_0_mult_485_C412_n344), .CI(dp_cluster_0_mult_485_C412_n358), 
        .CO(dp_cluster_0_mult_485_C412_n239), .S(
        dp_cluster_0_mult_485_C412_n240) );
  OAI22D1 U2073 ( .A1(n1967), .A2(n1970), .B1(n1966), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n373) );
  OAI22D1 U2074 ( .A1(n1951), .A2(n961), .B1(n1954), .B2(n1950), .ZN(
        dp_cluster_0_mult_485_C412_n358) );
  NR2D1 U2075 ( .A1(n1936), .A2(n1093), .ZN(dp_cluster_0_mult_485_C412_n344)
         );
  FA1D0 U2076 ( .A(dp_cluster_2_mult_485_C409_n373), .B(
        dp_cluster_2_mult_485_C409_n344), .CI(dp_cluster_2_mult_485_C409_n358), 
        .CO(dp_cluster_2_mult_485_C409_n239), .S(
        dp_cluster_2_mult_485_C409_n240) );
  OAI22D1 U2077 ( .A1(n2618), .A2(n2621), .B1(n2617), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n373) );
  OAI22D1 U2078 ( .A1(n2602), .A2(n985), .B1(n2605), .B2(n2601), .ZN(
        dp_cluster_2_mult_485_C409_n358) );
  NR2D1 U2079 ( .A1(n2587), .A2(n1090), .ZN(dp_cluster_2_mult_485_C409_n344)
         );
  FA1D0 U2080 ( .A(dp_cluster_1_mult_513_C418_n373), .B(
        dp_cluster_1_mult_513_C418_n344), .CI(dp_cluster_1_mult_513_C418_n358), 
        .CO(dp_cluster_1_mult_513_C418_n239), .S(
        dp_cluster_1_mult_513_C418_n240) );
  OAI22D1 U2081 ( .A1(n2141), .A2(n2144), .B1(n2140), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n373) );
  OAI22D1 U2082 ( .A1(n2125), .A2(n967), .B1(n2128), .B2(n2124), .ZN(
        dp_cluster_1_mult_513_C418_n358) );
  NR2D1 U2083 ( .A1(n2110), .A2(n1092), .ZN(dp_cluster_1_mult_513_C418_n344)
         );
  FA1D0 U2084 ( .A(dp_cluster_3_mult_513_C415_n373), .B(
        dp_cluster_3_mult_513_C415_n344), .CI(dp_cluster_3_mult_513_C415_n358), 
        .CO(dp_cluster_3_mult_513_C415_n239), .S(
        dp_cluster_3_mult_513_C415_n240) );
  OAI22D1 U2085 ( .A1(n2792), .A2(n2795), .B1(n2791), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n373) );
  OAI22D1 U2086 ( .A1(n2776), .A2(n991), .B1(n2779), .B2(n2775), .ZN(
        dp_cluster_3_mult_513_C415_n358) );
  NR2D1 U2087 ( .A1(n2761), .A2(n1089), .ZN(dp_cluster_3_mult_513_C415_n344)
         );
  FA1D0 U2088 ( .A(dp_cluster_1_mult_512_C418_n373), .B(
        dp_cluster_1_mult_512_C418_n344), .CI(dp_cluster_1_mult_512_C418_n358), 
        .CO(dp_cluster_1_mult_512_C418_n239), .S(
        dp_cluster_1_mult_512_C418_n240) );
  OAI22D1 U2089 ( .A1(n2293), .A2(n2296), .B1(n2292), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n373) );
  OAI22D1 U2090 ( .A1(n2277), .A2(n973), .B1(n2280), .B2(n2276), .ZN(
        dp_cluster_1_mult_512_C418_n358) );
  NR2D1 U2091 ( .A1(n2262), .A2(n1098), .ZN(dp_cluster_1_mult_512_C418_n344)
         );
  FA1D0 U2092 ( .A(dp_cluster_3_mult_512_C415_n373), .B(
        dp_cluster_3_mult_512_C415_n344), .CI(dp_cluster_3_mult_512_C415_n358), 
        .CO(dp_cluster_3_mult_512_C415_n239), .S(
        dp_cluster_3_mult_512_C415_n240) );
  OAI22D1 U2093 ( .A1(n2944), .A2(n2947), .B1(n2943), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n373) );
  OAI22D1 U2094 ( .A1(n2928), .A2(n997), .B1(n2931), .B2(n2927), .ZN(
        dp_cluster_3_mult_512_C415_n358) );
  NR2D1 U2095 ( .A1(n2913), .A2(n1095), .ZN(dp_cluster_3_mult_512_C415_n344)
         );
  FA1D0 U2096 ( .A(dp_cluster_0_mult_486_C412_n373), .B(
        dp_cluster_0_mult_486_C412_n344), .CI(dp_cluster_0_mult_486_C412_n358), 
        .CO(dp_cluster_0_mult_486_C412_n239), .S(
        dp_cluster_0_mult_486_C412_n240) );
  OAI22D1 U2097 ( .A1(n1815), .A2(n1818), .B1(n1814), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n373) );
  OAI22D1 U2098 ( .A1(n1799), .A2(n955), .B1(n1802), .B2(n1798), .ZN(
        dp_cluster_0_mult_486_C412_n358) );
  NR2D1 U2099 ( .A1(n1784), .A2(n1099), .ZN(dp_cluster_0_mult_486_C412_n344)
         );
  FA1D0 U2100 ( .A(dp_cluster_2_mult_486_C409_n373), .B(
        dp_cluster_2_mult_486_C409_n344), .CI(dp_cluster_2_mult_486_C409_n358), 
        .CO(dp_cluster_2_mult_486_C409_n239), .S(
        dp_cluster_2_mult_486_C409_n240) );
  OAI22D1 U2101 ( .A1(n2466), .A2(n2469), .B1(n2465), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n373) );
  OAI22D1 U2102 ( .A1(n2450), .A2(n979), .B1(n2453), .B2(n2449), .ZN(
        dp_cluster_2_mult_486_C409_n358) );
  NR2D1 U2103 ( .A1(n2435), .A2(n1096), .ZN(dp_cluster_2_mult_486_C409_n344)
         );
  OAI22D1 U2104 ( .A1(n1964), .A2(n1970), .B1(n1963), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n370) );
  OAI22D1 U2105 ( .A1(n1948), .A2(n961), .B1(n1954), .B2(n1947), .ZN(
        dp_cluster_0_mult_485_C412_n355) );
  OAI22D1 U2106 ( .A1(n1932), .A2(n960), .B1(n1936), .B2(n1931), .ZN(
        dp_cluster_0_mult_485_C412_n341) );
  OAI22D1 U2107 ( .A1(n2615), .A2(n2621), .B1(n2614), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n370) );
  OAI22D1 U2108 ( .A1(n2599), .A2(n985), .B1(n2605), .B2(n2598), .ZN(
        dp_cluster_2_mult_485_C409_n355) );
  OAI22D1 U2109 ( .A1(n2583), .A2(n984), .B1(n2587), .B2(n2582), .ZN(
        dp_cluster_2_mult_485_C409_n341) );
  OAI22D1 U2110 ( .A1(n2286), .A2(n2296), .B1(n2285), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n366) );
  OAI22D1 U2111 ( .A1(n2270), .A2(n973), .B1(n2280), .B2(n2269), .ZN(
        dp_cluster_1_mult_512_C418_n351) );
  OAI22D1 U2112 ( .A1(n2254), .A2(n972), .B1(n2262), .B2(n2253), .ZN(
        dp_cluster_1_mult_512_C418_n337) );
  OAI22D1 U2113 ( .A1(n2134), .A2(n2144), .B1(n2133), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n366) );
  OAI22D1 U2114 ( .A1(n2118), .A2(n967), .B1(n2128), .B2(n2117), .ZN(
        dp_cluster_1_mult_513_C418_n351) );
  OAI22D1 U2115 ( .A1(n2102), .A2(n966), .B1(n2110), .B2(n2101), .ZN(
        dp_cluster_1_mult_513_C418_n337) );
  OAI22D1 U2116 ( .A1(n1960), .A2(n1970), .B1(n1959), .B2(n1044), .ZN(
        dp_cluster_0_mult_485_C412_n366) );
  OAI22D1 U2117 ( .A1(n1944), .A2(n961), .B1(n1954), .B2(n1943), .ZN(
        dp_cluster_0_mult_485_C412_n351) );
  OAI22D1 U2118 ( .A1(n1928), .A2(n960), .B1(n1936), .B2(n1927), .ZN(
        dp_cluster_0_mult_485_C412_n337) );
  OAI22D1 U2119 ( .A1(n2937), .A2(n2947), .B1(n2936), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n366) );
  OAI22D1 U2120 ( .A1(n2921), .A2(n997), .B1(n2931), .B2(n2920), .ZN(
        dp_cluster_3_mult_512_C415_n351) );
  OAI22D1 U2121 ( .A1(n2905), .A2(n996), .B1(n2913), .B2(n2904), .ZN(
        dp_cluster_3_mult_512_C415_n337) );
  OAI22D1 U2122 ( .A1(n2785), .A2(n2795), .B1(n2784), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n366) );
  OAI22D1 U2123 ( .A1(n2769), .A2(n991), .B1(n2779), .B2(n2768), .ZN(
        dp_cluster_3_mult_513_C415_n351) );
  OAI22D1 U2124 ( .A1(n2753), .A2(n990), .B1(n2761), .B2(n2752), .ZN(
        dp_cluster_3_mult_513_C415_n337) );
  OAI22D1 U2125 ( .A1(n2611), .A2(n2621), .B1(n2610), .B2(n1022), .ZN(
        dp_cluster_2_mult_485_C409_n366) );
  OAI22D1 U2126 ( .A1(n2595), .A2(n985), .B1(n2605), .B2(n2594), .ZN(
        dp_cluster_2_mult_485_C409_n351) );
  OAI22D1 U2127 ( .A1(n2579), .A2(n984), .B1(n2587), .B2(n2578), .ZN(
        dp_cluster_2_mult_485_C409_n337) );
  OAI22D1 U2128 ( .A1(n1808), .A2(n1818), .B1(n1807), .B2(n1088), .ZN(
        dp_cluster_0_mult_486_C412_n366) );
  OAI22D1 U2129 ( .A1(n1792), .A2(n955), .B1(n1802), .B2(n1791), .ZN(
        dp_cluster_0_mult_486_C412_n351) );
  OAI22D1 U2130 ( .A1(n1776), .A2(n954), .B1(n1784), .B2(n1775), .ZN(
        dp_cluster_0_mult_486_C412_n337) );
  OAI22D1 U2131 ( .A1(n2459), .A2(n2469), .B1(n2458), .B2(n1066), .ZN(
        dp_cluster_2_mult_486_C409_n366) );
  OAI22D1 U2132 ( .A1(n2443), .A2(n979), .B1(n2453), .B2(n2442), .ZN(
        dp_cluster_2_mult_486_C409_n351) );
  OAI22D1 U2133 ( .A1(n2427), .A2(n978), .B1(n2435), .B2(n2426), .ZN(
        dp_cluster_2_mult_486_C409_n337) );
  OAI22D1 U2134 ( .A1(n2138), .A2(n2144), .B1(n2137), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n370) );
  OAI22D1 U2135 ( .A1(n2122), .A2(n967), .B1(n2128), .B2(n2121), .ZN(
        dp_cluster_1_mult_513_C418_n355) );
  OAI22D1 U2136 ( .A1(n2106), .A2(n966), .B1(n2110), .B2(n2105), .ZN(
        dp_cluster_1_mult_513_C418_n341) );
  OAI22D1 U2137 ( .A1(n2789), .A2(n2795), .B1(n2788), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n370) );
  OAI22D1 U2138 ( .A1(n2773), .A2(n991), .B1(n2779), .B2(n2772), .ZN(
        dp_cluster_3_mult_513_C415_n355) );
  OAI22D1 U2139 ( .A1(n2757), .A2(n990), .B1(n2761), .B2(n2756), .ZN(
        dp_cluster_3_mult_513_C415_n341) );
  OAI22D1 U2140 ( .A1(n2290), .A2(n2296), .B1(n2289), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n370) );
  OAI22D1 U2141 ( .A1(n2274), .A2(n973), .B1(n2280), .B2(n2273), .ZN(
        dp_cluster_1_mult_512_C418_n355) );
  OAI22D1 U2142 ( .A1(n2258), .A2(n972), .B1(n2262), .B2(n2257), .ZN(
        dp_cluster_1_mult_512_C418_n341) );
  OAI22D1 U2143 ( .A1(n1812), .A2(n1818), .B1(n1811), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n370) );
  OAI22D1 U2144 ( .A1(n1796), .A2(n955), .B1(n1802), .B2(n1795), .ZN(
        dp_cluster_0_mult_486_C412_n355) );
  OAI22D1 U2145 ( .A1(n1780), .A2(n954), .B1(n1784), .B2(n1779), .ZN(
        dp_cluster_0_mult_486_C412_n341) );
  OAI22D1 U2146 ( .A1(n2941), .A2(n2947), .B1(n2940), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n370) );
  OAI22D1 U2147 ( .A1(n2925), .A2(n997), .B1(n2931), .B2(n2924), .ZN(
        dp_cluster_3_mult_512_C415_n355) );
  OAI22D1 U2148 ( .A1(n2909), .A2(n996), .B1(n2913), .B2(n2908), .ZN(
        dp_cluster_3_mult_512_C415_n341) );
  OAI22D1 U2149 ( .A1(n2463), .A2(n2469), .B1(n2462), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n370) );
  OAI22D1 U2150 ( .A1(n2447), .A2(n979), .B1(n2453), .B2(n2446), .ZN(
        dp_cluster_2_mult_486_C409_n355) );
  OAI22D1 U2151 ( .A1(n2431), .A2(n978), .B1(n2435), .B2(n2430), .ZN(
        dp_cluster_2_mult_486_C409_n341) );
  FA1D0 U2152 ( .A(dp_cluster_0_mult_485_C412_n375), .B(
        dp_cluster_0_mult_485_C412_n360), .CI(dp_cluster_0_mult_485_C412_n77), 
        .CO(dp_cluster_0_mult_485_C412_n76), .S(dp_cluster_0_N59) );
  OAI22D1 U2153 ( .A1(n1969), .A2(n1970), .B1(n1968), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n375) );
  NR2D1 U2154 ( .A1(n1954), .A2(n1093), .ZN(dp_cluster_0_mult_485_C412_n360)
         );
  FA1D0 U2155 ( .A(dp_cluster_2_mult_485_C409_n375), .B(
        dp_cluster_2_mult_485_C409_n360), .CI(dp_cluster_2_mult_485_C409_n77), 
        .CO(dp_cluster_2_mult_485_C409_n76), .S(dp_cluster_2_N3) );
  OAI22D1 U2156 ( .A1(n2620), .A2(n2621), .B1(n2619), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n375) );
  NR2D1 U2157 ( .A1(n2605), .A2(n1090), .ZN(dp_cluster_2_mult_485_C409_n360)
         );
  FA1D0 U2158 ( .A(dp_cluster_0_mult_485_C412_n240), .B(
        dp_cluster_0_mult_485_C412_n241), .CI(dp_cluster_0_mult_485_C412_n75), 
        .CO(dp_cluster_0_mult_485_C412_n74), .S(dp_cluster_0_N61) );
  FA1D0 U2159 ( .A(dp_cluster_2_mult_485_C409_n240), .B(
        dp_cluster_2_mult_485_C409_n241), .CI(dp_cluster_2_mult_485_C409_n75), 
        .CO(dp_cluster_2_mult_485_C409_n74), .S(dp_cluster_2_N5) );
  OAI22D1 U2160 ( .A1(n2266), .A2(n973), .B1(n2280), .B2(n2265), .ZN(
        dp_cluster_1_mult_512_C418_n347) );
  OAI22D1 U2161 ( .A1(n2250), .A2(n972), .B1(n2262), .B2(n2249), .ZN(
        dp_cluster_1_mult_512_C418_n333) );
  OAI22D1 U2162 ( .A1(n2114), .A2(n967), .B1(n2128), .B2(n2113), .ZN(
        dp_cluster_1_mult_513_C418_n347) );
  OAI22D1 U2163 ( .A1(n2098), .A2(n966), .B1(n2110), .B2(n2097), .ZN(
        dp_cluster_1_mult_513_C418_n333) );
  OAI22D1 U2164 ( .A1(n1788), .A2(n955), .B1(n1802), .B2(n1787), .ZN(
        dp_cluster_0_mult_486_C412_n347) );
  OAI22D1 U2165 ( .A1(n1772), .A2(n954), .B1(n1784), .B2(n1771), .ZN(
        dp_cluster_0_mult_486_C412_n333) );
  OAI22D1 U2166 ( .A1(n1940), .A2(n961), .B1(n1954), .B2(n1939), .ZN(
        dp_cluster_0_mult_485_C412_n347) );
  OAI22D1 U2167 ( .A1(n1924), .A2(n960), .B1(n1936), .B2(n1923), .ZN(
        dp_cluster_0_mult_485_C412_n333) );
  OAI22D1 U2168 ( .A1(n2917), .A2(n997), .B1(n2931), .B2(n2916), .ZN(
        dp_cluster_3_mult_512_C415_n347) );
  OAI22D1 U2169 ( .A1(n2901), .A2(n996), .B1(n2913), .B2(n2900), .ZN(
        dp_cluster_3_mult_512_C415_n333) );
  OAI22D1 U2170 ( .A1(n2765), .A2(n991), .B1(n2779), .B2(n2764), .ZN(
        dp_cluster_3_mult_513_C415_n347) );
  OAI22D1 U2171 ( .A1(n2749), .A2(n990), .B1(n2761), .B2(n2748), .ZN(
        dp_cluster_3_mult_513_C415_n333) );
  OAI22D1 U2172 ( .A1(n2439), .A2(n979), .B1(n2453), .B2(n2438), .ZN(
        dp_cluster_2_mult_486_C409_n347) );
  OAI22D1 U2173 ( .A1(n2423), .A2(n978), .B1(n2435), .B2(n2422), .ZN(
        dp_cluster_2_mult_486_C409_n333) );
  OAI22D1 U2174 ( .A1(n2591), .A2(n985), .B1(n2605), .B2(n2590), .ZN(
        dp_cluster_2_mult_485_C409_n347) );
  OAI22D1 U2175 ( .A1(n2575), .A2(n984), .B1(n2587), .B2(n2574), .ZN(
        dp_cluster_2_mult_485_C409_n333) );
  IOA21D1 U2176 ( .A1(n1044), .A2(n2296), .B(n2281), .ZN(
        dp_cluster_1_mult_512_C418_n361) );
  OAI22D1 U2177 ( .A1(n2207), .A2(n971), .B1(n2300), .B2(n2206), .ZN(
        dp_cluster_1_mult_512_C418_n289) );
  OAI22D1 U2178 ( .A1(n2183), .A2(n2306), .B1(n2307), .B2(n2182), .ZN(
        dp_cluster_1_mult_512_C418_n262) );
  IOA21D1 U2179 ( .A1(n1088), .A2(n2144), .B(n2129), .ZN(
        dp_cluster_1_mult_513_C418_n361) );
  OAI22D1 U2180 ( .A1(n2055), .A2(n965), .B1(n2148), .B2(n2054), .ZN(
        dp_cluster_1_mult_513_C418_n289) );
  OAI22D1 U2181 ( .A1(n2031), .A2(n2154), .B1(n2155), .B2(n2030), .ZN(
        dp_cluster_1_mult_513_C418_n262) );
  IOA21D1 U2182 ( .A1(n1088), .A2(n1818), .B(n1803), .ZN(
        dp_cluster_0_mult_486_C412_n361) );
  OAI22D1 U2183 ( .A1(n1729), .A2(n953), .B1(n1822), .B2(n1728), .ZN(
        dp_cluster_0_mult_486_C412_n289) );
  OAI22D1 U2184 ( .A1(n1705), .A2(n1828), .B1(n1829), .B2(n1704), .ZN(
        dp_cluster_0_mult_486_C412_n262) );
  IOA21D1 U2185 ( .A1(n1044), .A2(n1970), .B(n1955), .ZN(
        dp_cluster_0_mult_485_C412_n361) );
  OAI22D1 U2186 ( .A1(n1881), .A2(n959), .B1(n1974), .B2(n1880), .ZN(
        dp_cluster_0_mult_485_C412_n289) );
  OAI22D1 U2187 ( .A1(n1857), .A2(n1980), .B1(n1981), .B2(n1856), .ZN(
        dp_cluster_0_mult_485_C412_n262) );
  IOA21D1 U2188 ( .A1(n1022), .A2(n2947), .B(n2932), .ZN(
        dp_cluster_3_mult_512_C415_n361) );
  OAI22D1 U2189 ( .A1(n2858), .A2(n995), .B1(n2951), .B2(n2857), .ZN(
        dp_cluster_3_mult_512_C415_n289) );
  OAI22D1 U2190 ( .A1(n2834), .A2(n2957), .B1(n2958), .B2(n2833), .ZN(
        dp_cluster_3_mult_512_C415_n262) );
  IOA21D1 U2191 ( .A1(n1066), .A2(n2795), .B(n2780), .ZN(
        dp_cluster_3_mult_513_C415_n361) );
  OAI22D1 U2192 ( .A1(n2706), .A2(n989), .B1(n2799), .B2(n2705), .ZN(
        dp_cluster_3_mult_513_C415_n289) );
  OAI22D1 U2193 ( .A1(n2682), .A2(n2805), .B1(n2806), .B2(n2681), .ZN(
        dp_cluster_3_mult_513_C415_n262) );
  IOA21D1 U2194 ( .A1(n1066), .A2(n2469), .B(n2454), .ZN(
        dp_cluster_2_mult_486_C409_n361) );
  OAI22D1 U2195 ( .A1(n2380), .A2(n977), .B1(n2473), .B2(n2379), .ZN(
        dp_cluster_2_mult_486_C409_n289) );
  OAI22D1 U2196 ( .A1(n2356), .A2(n2479), .B1(n2480), .B2(n2355), .ZN(
        dp_cluster_2_mult_486_C409_n262) );
  IOA21D1 U2197 ( .A1(n1022), .A2(n2621), .B(n2606), .ZN(
        dp_cluster_2_mult_485_C409_n361) );
  OAI22D1 U2198 ( .A1(n2532), .A2(n983), .B1(n2625), .B2(n2531), .ZN(
        dp_cluster_2_mult_485_C409_n289) );
  OAI22D1 U2199 ( .A1(n2508), .A2(n2631), .B1(n2632), .B2(n2507), .ZN(
        dp_cluster_2_mult_485_C409_n262) );
  XOR3D1 U2200 ( .A1(n2163), .A2(n2162), .A3(n2161), .Z(dp_cluster_1_N224) );
  XOR3D1 U2201 ( .A1(n2315), .A2(n2314), .A3(n2313), .Z(dp_cluster_1_N196) );
  OAI22D1 U2202 ( .A1(n2160), .A2(n969), .B1(n2158), .B2(n2157), .ZN(n2161) );
  XOR3D1 U2203 ( .A1(n2814), .A2(n2813), .A3(n2812), .Z(dp_cluster_3_N168) );
  XOR3D1 U2204 ( .A1(n2966), .A2(n2965), .A3(n2964), .Z(dp_cluster_3_N140) );
  OAI22D1 U2205 ( .A1(n2811), .A2(n993), .B1(n2809), .B2(n2808), .ZN(n2812) );
  OAI22D1 U2206 ( .A1(n1834), .A2(n957), .B1(n1832), .B2(n1831), .ZN(n1835) );
  OA22D0 U2207 ( .A1(n1830), .A2(n1829), .B1(n1828), .B2(n1827), .Z(n1837) );
  XOR3D1 U2208 ( .A1(dp_cluster_0_mult_486_C412_n81), .A2(
        dp_cluster_0_mult_486_C412_n80), .A3(dp_cluster_0_mult_486_C412_n52), 
        .Z(n1836) );
  OAI22D1 U2209 ( .A1(n2485), .A2(n981), .B1(n2483), .B2(n2482), .ZN(n2486) );
  OA22D0 U2210 ( .A1(n2481), .A2(n2480), .B1(n2479), .B2(n2478), .Z(n2488) );
  XOR3D1 U2211 ( .A1(dp_cluster_2_mult_486_C409_n81), .A2(
        dp_cluster_2_mult_486_C409_n80), .A3(dp_cluster_2_mult_486_C409_n52), 
        .Z(n2487) );
  FA1D0 U2212 ( .A(dp_cluster_0_mult_485_C412_n357), .B(
        dp_cluster_0_mult_485_C412_n372), .CI(dp_cluster_0_mult_485_C412_n238), 
        .CO(dp_cluster_0_mult_485_C412_n235), .S(
        dp_cluster_0_mult_485_C412_n236) );
  OAI22D1 U2213 ( .A1(n1966), .A2(n1970), .B1(n1965), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n372) );
  OAI22D1 U2214 ( .A1(n1950), .A2(n961), .B1(n1954), .B2(n1949), .ZN(
        dp_cluster_0_mult_485_C412_n357) );
  FA1D0 U2215 ( .A(dp_cluster_2_mult_485_C409_n357), .B(
        dp_cluster_2_mult_485_C409_n372), .CI(dp_cluster_2_mult_485_C409_n238), 
        .CO(dp_cluster_2_mult_485_C409_n235), .S(
        dp_cluster_2_mult_485_C409_n236) );
  OAI22D1 U2216 ( .A1(n2617), .A2(n2621), .B1(n2616), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n372) );
  OAI22D1 U2217 ( .A1(n2601), .A2(n985), .B1(n2605), .B2(n2600), .ZN(
        dp_cluster_2_mult_485_C409_n357) );
  FA1D0 U2218 ( .A(dp_cluster_1_mult_513_C418_n357), .B(
        dp_cluster_1_mult_513_C418_n372), .CI(dp_cluster_1_mult_513_C418_n238), 
        .CO(dp_cluster_1_mult_513_C418_n235), .S(
        dp_cluster_1_mult_513_C418_n236) );
  OAI22D1 U2219 ( .A1(n2140), .A2(n2144), .B1(n2139), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n372) );
  OAI22D1 U2220 ( .A1(n2124), .A2(n967), .B1(n2128), .B2(n2123), .ZN(
        dp_cluster_1_mult_513_C418_n357) );
  FA1D0 U2221 ( .A(dp_cluster_3_mult_513_C415_n357), .B(
        dp_cluster_3_mult_513_C415_n372), .CI(dp_cluster_3_mult_513_C415_n238), 
        .CO(dp_cluster_3_mult_513_C415_n235), .S(
        dp_cluster_3_mult_513_C415_n236) );
  OAI22D1 U2222 ( .A1(n2791), .A2(n2795), .B1(n2790), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n372) );
  OAI22D1 U2223 ( .A1(n2775), .A2(n991), .B1(n2779), .B2(n2774), .ZN(
        dp_cluster_3_mult_513_C415_n357) );
  FA1D0 U2224 ( .A(dp_cluster_1_mult_512_C418_n357), .B(
        dp_cluster_1_mult_512_C418_n372), .CI(dp_cluster_1_mult_512_C418_n238), 
        .CO(dp_cluster_1_mult_512_C418_n235), .S(
        dp_cluster_1_mult_512_C418_n236) );
  OAI22D1 U2225 ( .A1(n2292), .A2(n2296), .B1(n2291), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n372) );
  OAI22D1 U2226 ( .A1(n2276), .A2(n973), .B1(n2280), .B2(n2275), .ZN(
        dp_cluster_1_mult_512_C418_n357) );
  FA1D0 U2227 ( .A(dp_cluster_3_mult_512_C415_n357), .B(
        dp_cluster_3_mult_512_C415_n372), .CI(dp_cluster_3_mult_512_C415_n238), 
        .CO(dp_cluster_3_mult_512_C415_n235), .S(
        dp_cluster_3_mult_512_C415_n236) );
  OAI22D1 U2228 ( .A1(n2943), .A2(n2947), .B1(n2942), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n372) );
  OAI22D1 U2229 ( .A1(n2927), .A2(n997), .B1(n2931), .B2(n2926), .ZN(
        dp_cluster_3_mult_512_C415_n357) );
  FA1D0 U2230 ( .A(dp_cluster_0_mult_486_C412_n357), .B(
        dp_cluster_0_mult_486_C412_n372), .CI(dp_cluster_0_mult_486_C412_n238), 
        .CO(dp_cluster_0_mult_486_C412_n235), .S(
        dp_cluster_0_mult_486_C412_n236) );
  OAI22D1 U2231 ( .A1(n1814), .A2(n1818), .B1(n1813), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n372) );
  OAI22D1 U2232 ( .A1(n1798), .A2(n955), .B1(n1802), .B2(n1797), .ZN(
        dp_cluster_0_mult_486_C412_n357) );
  FA1D0 U2233 ( .A(dp_cluster_2_mult_486_C409_n357), .B(
        dp_cluster_2_mult_486_C409_n372), .CI(dp_cluster_2_mult_486_C409_n238), 
        .CO(dp_cluster_2_mult_486_C409_n235), .S(
        dp_cluster_2_mult_486_C409_n236) );
  OAI22D1 U2234 ( .A1(n2465), .A2(n2469), .B1(n2464), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n372) );
  OAI22D1 U2235 ( .A1(n2449), .A2(n979), .B1(n2453), .B2(n2448), .ZN(
        dp_cluster_2_mult_486_C409_n357) );
  CKBD1 U2236 ( .I(s1_7_r[2]), .Z(n1107) );
  CKBD1 U2237 ( .I(s1_5_r[2]), .Z(n1110) );
  CKBD1 U2238 ( .I(s1_7_i[2]), .Z(n1101) );
  CKBD1 U2239 ( .I(s1_5_i[2]), .Z(n1104) );
  FA1D0 U2240 ( .A(dp_cluster_1_mult_513_C418_n240), .B(
        dp_cluster_1_mult_513_C418_n241), .CI(dp_cluster_1_mult_513_C418_n75), 
        .CO(dp_cluster_1_mult_513_C418_n74), .S(dp_cluster_1_N201) );
  FA1D0 U2241 ( .A(dp_cluster_3_mult_513_C415_n240), .B(
        dp_cluster_3_mult_513_C415_n241), .CI(dp_cluster_3_mult_513_C415_n75), 
        .CO(dp_cluster_3_mult_513_C415_n74), .S(dp_cluster_3_N145) );
  FA1D0 U2242 ( .A(dp_cluster_1_mult_512_C418_n240), .B(
        dp_cluster_1_mult_512_C418_n241), .CI(dp_cluster_1_mult_512_C418_n75), 
        .CO(dp_cluster_1_mult_512_C418_n74), .S(dp_cluster_1_N173) );
  FA1D0 U2243 ( .A(dp_cluster_3_mult_512_C415_n240), .B(
        dp_cluster_3_mult_512_C415_n241), .CI(dp_cluster_3_mult_512_C415_n75), 
        .CO(dp_cluster_3_mult_512_C415_n74), .S(dp_cluster_3_N117) );
  FA1D0 U2244 ( .A(dp_cluster_1_mult_513_C418_n375), .B(
        dp_cluster_1_mult_513_C418_n360), .CI(dp_cluster_1_mult_513_C418_n77), 
        .CO(dp_cluster_1_mult_513_C418_n76), .S(dp_cluster_1_N199) );
  OAI22D1 U2245 ( .A1(n2143), .A2(n2144), .B1(n2142), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n375) );
  NR2D1 U2246 ( .A1(n2128), .A2(n1092), .ZN(dp_cluster_1_mult_513_C418_n360)
         );
  FA1D0 U2247 ( .A(dp_cluster_3_mult_513_C415_n375), .B(
        dp_cluster_3_mult_513_C415_n360), .CI(dp_cluster_3_mult_513_C415_n77), 
        .CO(dp_cluster_3_mult_513_C415_n76), .S(dp_cluster_3_N143) );
  OAI22D1 U2248 ( .A1(n2794), .A2(n2795), .B1(n2793), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n375) );
  NR2D1 U2249 ( .A1(n2779), .A2(n1089), .ZN(dp_cluster_3_mult_513_C415_n360)
         );
  FA1D0 U2250 ( .A(dp_cluster_1_mult_512_C418_n375), .B(
        dp_cluster_1_mult_512_C418_n360), .CI(dp_cluster_1_mult_512_C418_n77), 
        .CO(dp_cluster_1_mult_512_C418_n76), .S(dp_cluster_1_N171) );
  OAI22D1 U2251 ( .A1(n2295), .A2(n2296), .B1(n2294), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n375) );
  NR2D1 U2252 ( .A1(n2280), .A2(n1098), .ZN(dp_cluster_1_mult_512_C418_n360)
         );
  FA1D0 U2253 ( .A(dp_cluster_3_mult_512_C415_n375), .B(
        dp_cluster_3_mult_512_C415_n360), .CI(dp_cluster_3_mult_512_C415_n77), 
        .CO(dp_cluster_3_mult_512_C415_n76), .S(dp_cluster_3_N115) );
  OAI22D1 U2254 ( .A1(n2946), .A2(n2947), .B1(n2945), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n375) );
  NR2D1 U2255 ( .A1(n2931), .A2(n1095), .ZN(dp_cluster_3_mult_512_C415_n360)
         );
  HA1D0 U2256 ( .A(dp_cluster_0_mult_485_C412_n359), .B(
        dp_cluster_0_mult_485_C412_n374), .CO(dp_cluster_0_mult_485_C412_n241), 
        .S(dp_cluster_0_mult_485_C412_n242) );
  OAI22D1 U2257 ( .A1(n1968), .A2(n1970), .B1(n1967), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n374) );
  OAI22D1 U2258 ( .A1(n1953), .A2(n961), .B1(n1954), .B2(n1951), .ZN(
        dp_cluster_0_mult_485_C412_n359) );
  HA1D0 U2259 ( .A(dp_cluster_2_mult_485_C409_n359), .B(
        dp_cluster_2_mult_485_C409_n374), .CO(dp_cluster_2_mult_485_C409_n241), 
        .S(dp_cluster_2_mult_485_C409_n242) );
  OAI22D1 U2260 ( .A1(n2619), .A2(n2621), .B1(n2618), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n374) );
  OAI22D1 U2261 ( .A1(n2604), .A2(n985), .B1(n2605), .B2(n2602), .ZN(
        dp_cluster_2_mult_485_C409_n359) );
  HA1D0 U2262 ( .A(dp_cluster_1_mult_513_C418_n359), .B(
        dp_cluster_1_mult_513_C418_n374), .CO(dp_cluster_1_mult_513_C418_n241), 
        .S(dp_cluster_1_mult_513_C418_n242) );
  OAI22D1 U2263 ( .A1(n2142), .A2(n2144), .B1(n2141), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n374) );
  OAI22D1 U2264 ( .A1(n2127), .A2(n967), .B1(n2128), .B2(n2125), .ZN(
        dp_cluster_1_mult_513_C418_n359) );
  HA1D0 U2265 ( .A(dp_cluster_3_mult_513_C415_n359), .B(
        dp_cluster_3_mult_513_C415_n374), .CO(dp_cluster_3_mult_513_C415_n241), 
        .S(dp_cluster_3_mult_513_C415_n242) );
  OAI22D1 U2266 ( .A1(n2793), .A2(n2795), .B1(n2792), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n374) );
  OAI22D1 U2267 ( .A1(n2778), .A2(n991), .B1(n2779), .B2(n2776), .ZN(
        dp_cluster_3_mult_513_C415_n359) );
  HA1D0 U2268 ( .A(dp_cluster_1_mult_512_C418_n359), .B(
        dp_cluster_1_mult_512_C418_n374), .CO(dp_cluster_1_mult_512_C418_n241), 
        .S(dp_cluster_1_mult_512_C418_n242) );
  OAI22D1 U2269 ( .A1(n2294), .A2(n2296), .B1(n2293), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n374) );
  OAI22D1 U2270 ( .A1(n2279), .A2(n973), .B1(n2280), .B2(n2277), .ZN(
        dp_cluster_1_mult_512_C418_n359) );
  HA1D0 U2271 ( .A(dp_cluster_3_mult_512_C415_n359), .B(
        dp_cluster_3_mult_512_C415_n374), .CO(dp_cluster_3_mult_512_C415_n241), 
        .S(dp_cluster_3_mult_512_C415_n242) );
  OAI22D1 U2272 ( .A1(n2945), .A2(n2947), .B1(n2944), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n374) );
  OAI22D1 U2273 ( .A1(n2930), .A2(n997), .B1(n2931), .B2(n2928), .ZN(
        dp_cluster_3_mult_512_C415_n359) );
  HA1D0 U2274 ( .A(dp_cluster_0_mult_486_C412_n359), .B(
        dp_cluster_0_mult_486_C412_n374), .CO(dp_cluster_0_mult_486_C412_n241), 
        .S(dp_cluster_0_mult_486_C412_n242) );
  OAI22D1 U2275 ( .A1(n1816), .A2(n1818), .B1(n1815), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n374) );
  OAI22D1 U2276 ( .A1(n1801), .A2(n955), .B1(n1802), .B2(n1799), .ZN(
        dp_cluster_0_mult_486_C412_n359) );
  HA1D0 U2277 ( .A(dp_cluster_2_mult_486_C409_n359), .B(
        dp_cluster_2_mult_486_C409_n374), .CO(dp_cluster_2_mult_486_C409_n241), 
        .S(dp_cluster_2_mult_486_C409_n242) );
  OAI22D1 U2278 ( .A1(n2467), .A2(n2469), .B1(n2466), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n374) );
  OAI22D1 U2279 ( .A1(n2452), .A2(n979), .B1(n2453), .B2(n2450), .ZN(
        dp_cluster_2_mult_486_C409_n359) );
  OAI22D1 U2280 ( .A1(n2285), .A2(n2296), .B1(n2284), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n365) );
  OAI22D1 U2281 ( .A1(n2269), .A2(n973), .B1(n2280), .B2(n2268), .ZN(
        dp_cluster_1_mult_512_C418_n350) );
  OAI22D1 U2282 ( .A1(n2237), .A2(n974), .B1(n2244), .B2(n2236), .ZN(
        dp_cluster_1_mult_512_C418_n322) );
  OAI22D1 U2283 ( .A1(n2133), .A2(n2144), .B1(n2132), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n365) );
  OAI22D1 U2284 ( .A1(n2117), .A2(n967), .B1(n2128), .B2(n2116), .ZN(
        dp_cluster_1_mult_513_C418_n350) );
  OAI22D1 U2285 ( .A1(n2085), .A2(n968), .B1(n2092), .B2(n2084), .ZN(
        dp_cluster_1_mult_513_C418_n322) );
  OAI22D1 U2286 ( .A1(n1807), .A2(n1818), .B1(n1806), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n365) );
  OAI22D1 U2287 ( .A1(n1791), .A2(n955), .B1(n1802), .B2(n1790), .ZN(
        dp_cluster_0_mult_486_C412_n350) );
  OAI22D1 U2288 ( .A1(n1759), .A2(n956), .B1(n1766), .B2(n1758), .ZN(
        dp_cluster_0_mult_486_C412_n322) );
  OAI22D1 U2289 ( .A1(n1959), .A2(n1970), .B1(n1958), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n365) );
  OAI22D1 U2290 ( .A1(n1943), .A2(n961), .B1(n1954), .B2(n1942), .ZN(
        dp_cluster_0_mult_485_C412_n350) );
  OAI22D1 U2291 ( .A1(n1911), .A2(n962), .B1(n1918), .B2(n1910), .ZN(
        dp_cluster_0_mult_485_C412_n322) );
  OAI22D1 U2292 ( .A1(n2936), .A2(n2947), .B1(n2935), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n365) );
  OAI22D1 U2293 ( .A1(n2920), .A2(n997), .B1(n2931), .B2(n2919), .ZN(
        dp_cluster_3_mult_512_C415_n350) );
  OAI22D1 U2294 ( .A1(n2888), .A2(n998), .B1(n2895), .B2(n2887), .ZN(
        dp_cluster_3_mult_512_C415_n322) );
  OAI22D1 U2295 ( .A1(n2784), .A2(n2795), .B1(n2783), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n365) );
  OAI22D1 U2296 ( .A1(n2768), .A2(n991), .B1(n2779), .B2(n2767), .ZN(
        dp_cluster_3_mult_513_C415_n350) );
  OAI22D1 U2297 ( .A1(n2736), .A2(n992), .B1(n2743), .B2(n2735), .ZN(
        dp_cluster_3_mult_513_C415_n322) );
  OAI22D1 U2298 ( .A1(n2458), .A2(n2469), .B1(n2457), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n365) );
  OAI22D1 U2299 ( .A1(n2442), .A2(n979), .B1(n2453), .B2(n2441), .ZN(
        dp_cluster_2_mult_486_C409_n350) );
  OAI22D1 U2300 ( .A1(n2410), .A2(n980), .B1(n2417), .B2(n2409), .ZN(
        dp_cluster_2_mult_486_C409_n322) );
  OAI22D1 U2301 ( .A1(n2610), .A2(n2621), .B1(n2609), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n365) );
  OAI22D1 U2302 ( .A1(n2594), .A2(n985), .B1(n2605), .B2(n2593), .ZN(
        dp_cluster_2_mult_485_C409_n350) );
  OAI22D1 U2303 ( .A1(n2562), .A2(n986), .B1(n2569), .B2(n2561), .ZN(
        dp_cluster_2_mult_485_C409_n322) );
  OAI22D1 U2304 ( .A1(n2268), .A2(n973), .B1(n2280), .B2(n2267), .ZN(
        dp_cluster_1_mult_512_C418_n349) );
  OAI22D1 U2305 ( .A1(n2252), .A2(n972), .B1(n2262), .B2(n2251), .ZN(
        dp_cluster_1_mult_512_C418_n335) );
  OAI22D1 U2306 ( .A1(n2222), .A2(n976), .B1(n2304), .B2(n2221), .ZN(
        dp_cluster_1_mult_512_C418_n306) );
  OAI22D1 U2307 ( .A1(n2116), .A2(n967), .B1(n2128), .B2(n2115), .ZN(
        dp_cluster_1_mult_513_C418_n349) );
  OAI22D1 U2308 ( .A1(n2100), .A2(n966), .B1(n2110), .B2(n2099), .ZN(
        dp_cluster_1_mult_513_C418_n335) );
  OAI22D1 U2309 ( .A1(n2070), .A2(n970), .B1(n2152), .B2(n2069), .ZN(
        dp_cluster_1_mult_513_C418_n306) );
  OAI22D1 U2310 ( .A1(n1790), .A2(n955), .B1(n1802), .B2(n1789), .ZN(
        dp_cluster_0_mult_486_C412_n349) );
  OAI22D1 U2311 ( .A1(n1774), .A2(n954), .B1(n1784), .B2(n1773), .ZN(
        dp_cluster_0_mult_486_C412_n335) );
  OAI22D1 U2312 ( .A1(n1744), .A2(n958), .B1(n1826), .B2(n1743), .ZN(
        dp_cluster_0_mult_486_C412_n306) );
  OAI22D1 U2313 ( .A1(n1942), .A2(n961), .B1(n1954), .B2(n1941), .ZN(
        dp_cluster_0_mult_485_C412_n349) );
  OAI22D1 U2314 ( .A1(n1926), .A2(n960), .B1(n1936), .B2(n1925), .ZN(
        dp_cluster_0_mult_485_C412_n335) );
  OAI22D1 U2315 ( .A1(n1896), .A2(n964), .B1(n1978), .B2(n1895), .ZN(
        dp_cluster_0_mult_485_C412_n306) );
  OAI22D1 U2316 ( .A1(n2919), .A2(n997), .B1(n2931), .B2(n2918), .ZN(
        dp_cluster_3_mult_512_C415_n349) );
  OAI22D1 U2317 ( .A1(n2903), .A2(n996), .B1(n2913), .B2(n2902), .ZN(
        dp_cluster_3_mult_512_C415_n335) );
  OAI22D1 U2318 ( .A1(n2873), .A2(n1000), .B1(n2955), .B2(n2872), .ZN(
        dp_cluster_3_mult_512_C415_n306) );
  OAI22D1 U2319 ( .A1(n2767), .A2(n991), .B1(n2779), .B2(n2766), .ZN(
        dp_cluster_3_mult_513_C415_n349) );
  OAI22D1 U2320 ( .A1(n2751), .A2(n990), .B1(n2761), .B2(n2750), .ZN(
        dp_cluster_3_mult_513_C415_n335) );
  OAI22D1 U2321 ( .A1(n2721), .A2(n994), .B1(n2803), .B2(n2720), .ZN(
        dp_cluster_3_mult_513_C415_n306) );
  OAI22D1 U2322 ( .A1(n2441), .A2(n979), .B1(n2453), .B2(n2440), .ZN(
        dp_cluster_2_mult_486_C409_n349) );
  OAI22D1 U2323 ( .A1(n2425), .A2(n978), .B1(n2435), .B2(n2424), .ZN(
        dp_cluster_2_mult_486_C409_n335) );
  OAI22D1 U2324 ( .A1(n2395), .A2(n982), .B1(n2477), .B2(n2394), .ZN(
        dp_cluster_2_mult_486_C409_n306) );
  OAI22D1 U2325 ( .A1(n2593), .A2(n985), .B1(n2605), .B2(n2592), .ZN(
        dp_cluster_2_mult_485_C409_n349) );
  OAI22D1 U2326 ( .A1(n2577), .A2(n984), .B1(n2587), .B2(n2576), .ZN(
        dp_cluster_2_mult_485_C409_n335) );
  OAI22D1 U2327 ( .A1(n2547), .A2(n988), .B1(n2629), .B2(n2546), .ZN(
        dp_cluster_2_mult_485_C409_n306) );
  OAI22D1 U2328 ( .A1(n2283), .A2(n2296), .B1(n2282), .B2(n1043), .ZN(
        dp_cluster_1_mult_512_C418_n363) );
  OAI22D1 U2329 ( .A1(n2267), .A2(n973), .B1(n2280), .B2(n2266), .ZN(
        dp_cluster_1_mult_512_C418_n348) );
  OAI22D1 U2330 ( .A1(n2251), .A2(n972), .B1(n2262), .B2(n2250), .ZN(
        dp_cluster_1_mult_512_C418_n334) );
  OAI22D1 U2331 ( .A1(n2131), .A2(n2144), .B1(n2130), .B2(n1087), .ZN(
        dp_cluster_1_mult_513_C418_n363) );
  OAI22D1 U2332 ( .A1(n2115), .A2(n967), .B1(n2128), .B2(n2114), .ZN(
        dp_cluster_1_mult_513_C418_n348) );
  OAI22D1 U2333 ( .A1(n2099), .A2(n966), .B1(n2110), .B2(n2098), .ZN(
        dp_cluster_1_mult_513_C418_n334) );
  OAI22D1 U2334 ( .A1(n1805), .A2(n1818), .B1(n1804), .B2(n1088), .ZN(
        dp_cluster_0_mult_486_C412_n363) );
  OAI22D1 U2335 ( .A1(n1789), .A2(n955), .B1(n1802), .B2(n1788), .ZN(
        dp_cluster_0_mult_486_C412_n348) );
  OAI22D1 U2336 ( .A1(n1773), .A2(n954), .B1(n1784), .B2(n1772), .ZN(
        dp_cluster_0_mult_486_C412_n334) );
  OAI22D1 U2337 ( .A1(n1957), .A2(n1970), .B1(n1956), .B2(n1044), .ZN(
        dp_cluster_0_mult_485_C412_n363) );
  OAI22D1 U2338 ( .A1(n1941), .A2(n961), .B1(n1954), .B2(n1940), .ZN(
        dp_cluster_0_mult_485_C412_n348) );
  OAI22D1 U2339 ( .A1(n1925), .A2(n960), .B1(n1936), .B2(n1924), .ZN(
        dp_cluster_0_mult_485_C412_n334) );
  OAI22D1 U2340 ( .A1(n2934), .A2(n2947), .B1(n2933), .B2(n1021), .ZN(
        dp_cluster_3_mult_512_C415_n363) );
  OAI22D1 U2341 ( .A1(n2918), .A2(n997), .B1(n2931), .B2(n2917), .ZN(
        dp_cluster_3_mult_512_C415_n348) );
  OAI22D1 U2342 ( .A1(n2902), .A2(n996), .B1(n2913), .B2(n2901), .ZN(
        dp_cluster_3_mult_512_C415_n334) );
  OAI22D1 U2343 ( .A1(n2782), .A2(n2795), .B1(n2781), .B2(n1065), .ZN(
        dp_cluster_3_mult_513_C415_n363) );
  OAI22D1 U2344 ( .A1(n2766), .A2(n991), .B1(n2779), .B2(n2765), .ZN(
        dp_cluster_3_mult_513_C415_n348) );
  OAI22D1 U2345 ( .A1(n2750), .A2(n990), .B1(n2761), .B2(n2749), .ZN(
        dp_cluster_3_mult_513_C415_n334) );
  OAI22D1 U2346 ( .A1(n2456), .A2(n2469), .B1(n2455), .B2(n1066), .ZN(
        dp_cluster_2_mult_486_C409_n363) );
  OAI22D1 U2347 ( .A1(n2440), .A2(n979), .B1(n2453), .B2(n2439), .ZN(
        dp_cluster_2_mult_486_C409_n348) );
  OAI22D1 U2348 ( .A1(n2424), .A2(n978), .B1(n2435), .B2(n2423), .ZN(
        dp_cluster_2_mult_486_C409_n334) );
  OAI22D1 U2349 ( .A1(n2608), .A2(n2621), .B1(n2607), .B2(n1022), .ZN(
        dp_cluster_2_mult_485_C409_n363) );
  OAI22D1 U2350 ( .A1(n2592), .A2(n985), .B1(n2605), .B2(n2591), .ZN(
        dp_cluster_2_mult_485_C409_n348) );
  OAI22D1 U2351 ( .A1(n2576), .A2(n984), .B1(n2587), .B2(n2575), .ZN(
        dp_cluster_2_mult_485_C409_n334) );
  OAI22D1 U2352 ( .A1(n2228), .A2(n974), .B1(n2244), .B2(n2227), .ZN(
        dp_cluster_1_mult_512_C418_n313) );
  OAI22D1 U2353 ( .A1(n2214), .A2(n976), .B1(n2304), .B2(n2213), .ZN(
        dp_cluster_1_mult_512_C418_n298) );
  INVD1 U2354 ( .I(dp_cluster_1_mult_512_C418_n112), .ZN(n1157) );
  OAI22D1 U2355 ( .A1(n2076), .A2(n968), .B1(n2092), .B2(n2075), .ZN(
        dp_cluster_1_mult_513_C418_n313) );
  OAI22D1 U2356 ( .A1(n2062), .A2(n970), .B1(n2152), .B2(n2061), .ZN(
        dp_cluster_1_mult_513_C418_n298) );
  INVD1 U2357 ( .I(dp_cluster_1_mult_513_C418_n112), .ZN(n1292) );
  OAI22D1 U2358 ( .A1(n1750), .A2(n956), .B1(n1766), .B2(n1749), .ZN(
        dp_cluster_0_mult_486_C412_n313) );
  OAI22D1 U2359 ( .A1(n1736), .A2(n958), .B1(n1826), .B2(n1735), .ZN(
        dp_cluster_0_mult_486_C412_n298) );
  INVD1 U2360 ( .I(dp_cluster_0_mult_486_C412_n112), .ZN(n1290) );
  OAI22D1 U2361 ( .A1(n1902), .A2(n962), .B1(n1918), .B2(n1901), .ZN(
        dp_cluster_0_mult_485_C412_n313) );
  OAI22D1 U2362 ( .A1(n1888), .A2(n964), .B1(n1978), .B2(n1887), .ZN(
        dp_cluster_0_mult_485_C412_n298) );
  INVD1 U2363 ( .I(dp_cluster_0_mult_485_C412_n112), .ZN(n1154) );
  OAI22D1 U2364 ( .A1(n2879), .A2(n998), .B1(n2895), .B2(n2878), .ZN(
        dp_cluster_3_mult_512_C415_n313) );
  OAI22D1 U2365 ( .A1(n2865), .A2(n1000), .B1(n2955), .B2(n2864), .ZN(
        dp_cluster_3_mult_512_C415_n298) );
  INVD1 U2366 ( .I(dp_cluster_3_mult_512_C415_n112), .ZN(n1118) );
  OAI22D1 U2367 ( .A1(n2727), .A2(n992), .B1(n2743), .B2(n2726), .ZN(
        dp_cluster_3_mult_513_C415_n313) );
  OAI22D1 U2368 ( .A1(n2713), .A2(n994), .B1(n2803), .B2(n2712), .ZN(
        dp_cluster_3_mult_513_C415_n298) );
  INVD1 U2369 ( .I(dp_cluster_3_mult_513_C415_n112), .ZN(n1259) );
  OAI22D1 U2370 ( .A1(n2401), .A2(n980), .B1(n2417), .B2(n2400), .ZN(
        dp_cluster_2_mult_486_C409_n313) );
  OAI22D1 U2371 ( .A1(n2387), .A2(n982), .B1(n2477), .B2(n2386), .ZN(
        dp_cluster_2_mult_486_C409_n298) );
  INVD1 U2372 ( .I(dp_cluster_2_mult_486_C409_n112), .ZN(n1257) );
  OAI22D1 U2373 ( .A1(n2553), .A2(n986), .B1(n2569), .B2(n2552), .ZN(
        dp_cluster_2_mult_485_C409_n313) );
  OAI22D1 U2374 ( .A1(n2539), .A2(n988), .B1(n2629), .B2(n2538), .ZN(
        dp_cluster_2_mult_485_C409_n298) );
  INVD1 U2375 ( .I(dp_cluster_2_mult_485_C409_n112), .ZN(n1115) );
  OAI22D1 U2376 ( .A1(n2213), .A2(n976), .B1(n2304), .B2(n2302), .ZN(
        dp_cluster_1_mult_512_C418_n297) );
  OAI22D1 U2377 ( .A1(n2201), .A2(n971), .B1(n2300), .B2(n2200), .ZN(
        dp_cluster_1_mult_512_C418_n284) );
  OAI22D1 U2378 ( .A1(n2061), .A2(n970), .B1(n2152), .B2(n2150), .ZN(
        dp_cluster_1_mult_513_C418_n297) );
  OAI22D1 U2379 ( .A1(n2049), .A2(n965), .B1(n2148), .B2(n2048), .ZN(
        dp_cluster_1_mult_513_C418_n284) );
  OAI22D1 U2380 ( .A1(n1735), .A2(n958), .B1(n1826), .B2(n1824), .ZN(
        dp_cluster_0_mult_486_C412_n297) );
  OAI22D1 U2381 ( .A1(n1723), .A2(n953), .B1(n1822), .B2(n1722), .ZN(
        dp_cluster_0_mult_486_C412_n284) );
  OAI22D1 U2382 ( .A1(n1887), .A2(n964), .B1(n1978), .B2(n1976), .ZN(
        dp_cluster_0_mult_485_C412_n297) );
  OAI22D1 U2383 ( .A1(n1875), .A2(n959), .B1(n1974), .B2(n1874), .ZN(
        dp_cluster_0_mult_485_C412_n284) );
  OAI22D1 U2384 ( .A1(n2864), .A2(n1000), .B1(n2955), .B2(n2953), .ZN(
        dp_cluster_3_mult_512_C415_n297) );
  OAI22D1 U2385 ( .A1(n2852), .A2(n995), .B1(n2951), .B2(n2851), .ZN(
        dp_cluster_3_mult_512_C415_n284) );
  OAI22D1 U2386 ( .A1(n2712), .A2(n994), .B1(n2803), .B2(n2801), .ZN(
        dp_cluster_3_mult_513_C415_n297) );
  OAI22D1 U2387 ( .A1(n2700), .A2(n989), .B1(n2799), .B2(n2699), .ZN(
        dp_cluster_3_mult_513_C415_n284) );
  OAI22D1 U2388 ( .A1(n2386), .A2(n982), .B1(n2477), .B2(n2475), .ZN(
        dp_cluster_2_mult_486_C409_n297) );
  OAI22D1 U2389 ( .A1(n2374), .A2(n977), .B1(n2473), .B2(n2373), .ZN(
        dp_cluster_2_mult_486_C409_n284) );
  OAI22D1 U2390 ( .A1(n2538), .A2(n988), .B1(n2629), .B2(n2627), .ZN(
        dp_cluster_2_mult_485_C409_n297) );
  OAI22D1 U2391 ( .A1(n2526), .A2(n983), .B1(n2625), .B2(n2525), .ZN(
        dp_cluster_2_mult_485_C409_n284) );
  OAI22D1 U2392 ( .A1(n2255), .A2(n972), .B1(n2262), .B2(n2254), .ZN(
        dp_cluster_1_mult_512_C418_n338) );
  OAI22D1 U2393 ( .A1(n2239), .A2(n974), .B1(n2244), .B2(n2238), .ZN(
        dp_cluster_1_mult_512_C418_n324) );
  NR2D1 U2394 ( .A1(n2300), .A2(n1098), .ZN(dp_cluster_1_mult_512_C418_n295)
         );
  OAI22D1 U2395 ( .A1(n2103), .A2(n966), .B1(n2110), .B2(n2102), .ZN(
        dp_cluster_1_mult_513_C418_n338) );
  OAI22D1 U2396 ( .A1(n2087), .A2(n968), .B1(n2092), .B2(n2086), .ZN(
        dp_cluster_1_mult_513_C418_n324) );
  NR2D1 U2397 ( .A1(n2148), .A2(n1092), .ZN(dp_cluster_1_mult_513_C418_n295)
         );
  OAI22D1 U2398 ( .A1(n1929), .A2(n960), .B1(n1936), .B2(n1928), .ZN(
        dp_cluster_0_mult_485_C412_n338) );
  OAI22D1 U2399 ( .A1(n1913), .A2(n962), .B1(n1918), .B2(n1912), .ZN(
        dp_cluster_0_mult_485_C412_n324) );
  NR2D1 U2400 ( .A1(n1974), .A2(n1093), .ZN(dp_cluster_0_mult_485_C412_n295)
         );
  OAI22D1 U2401 ( .A1(n2906), .A2(n996), .B1(n2913), .B2(n2905), .ZN(
        dp_cluster_3_mult_512_C415_n338) );
  OAI22D1 U2402 ( .A1(n2890), .A2(n998), .B1(n2895), .B2(n2889), .ZN(
        dp_cluster_3_mult_512_C415_n324) );
  NR2D1 U2403 ( .A1(n2951), .A2(n1095), .ZN(dp_cluster_3_mult_512_C415_n295)
         );
  OAI22D1 U2404 ( .A1(n2754), .A2(n990), .B1(n2761), .B2(n2753), .ZN(
        dp_cluster_3_mult_513_C415_n338) );
  OAI22D1 U2405 ( .A1(n2738), .A2(n992), .B1(n2743), .B2(n2737), .ZN(
        dp_cluster_3_mult_513_C415_n324) );
  NR2D1 U2406 ( .A1(n2799), .A2(n1089), .ZN(dp_cluster_3_mult_513_C415_n295)
         );
  OAI22D1 U2407 ( .A1(n2580), .A2(n984), .B1(n2587), .B2(n2579), .ZN(
        dp_cluster_2_mult_485_C409_n338) );
  OAI22D1 U2408 ( .A1(n2564), .A2(n986), .B1(n2569), .B2(n2563), .ZN(
        dp_cluster_2_mult_485_C409_n324) );
  NR2D1 U2409 ( .A1(n2625), .A2(n1090), .ZN(dp_cluster_2_mult_485_C409_n295)
         );
  OAI22D1 U2410 ( .A1(n1777), .A2(n954), .B1(n1784), .B2(n1776), .ZN(
        dp_cluster_0_mult_486_C412_n338) );
  OAI22D1 U2411 ( .A1(n1761), .A2(n956), .B1(n1766), .B2(n1760), .ZN(
        dp_cluster_0_mult_486_C412_n324) );
  NR2D1 U2412 ( .A1(n1822), .A2(n1099), .ZN(dp_cluster_0_mult_486_C412_n295)
         );
  OAI22D1 U2413 ( .A1(n2428), .A2(n978), .B1(n2435), .B2(n2427), .ZN(
        dp_cluster_2_mult_486_C409_n338) );
  OAI22D1 U2414 ( .A1(n2412), .A2(n980), .B1(n2417), .B2(n2411), .ZN(
        dp_cluster_2_mult_486_C409_n324) );
  NR2D1 U2415 ( .A1(n2473), .A2(n1096), .ZN(dp_cluster_2_mult_486_C409_n295)
         );
  CKBD1 U2416 ( .I(n1952), .Z(n961) );
  ND2D1 U2417 ( .A1(n1954), .A2(n1840), .ZN(n1952) );
  CKBD1 U2418 ( .I(n2603), .Z(n985) );
  ND2D1 U2419 ( .A1(n2605), .A2(n2491), .ZN(n2603) );
  CKBD1 U2420 ( .I(n1800), .Z(n955) );
  ND2D1 U2421 ( .A1(n1802), .A2(n1688), .ZN(n1800) );
  CKBD1 U2422 ( .I(n2451), .Z(n979) );
  ND2D1 U2423 ( .A1(n2453), .A2(n2339), .ZN(n2451) );
  IOA21D1 U2424 ( .A1(n2320), .A2(dp_cluster_1_N172), .B(n2319), .ZN(n2322) );
  OAI21D1 U2425 ( .A1(dp_cluster_1_N172), .A2(n2320), .B(dp_cluster_1_N200), 
        .ZN(n2319) );
  IOA21D1 U2426 ( .A1(n2318), .A2(dp_cluster_1_N171), .B(n2317), .ZN(n2320) );
  OAI21D1 U2427 ( .A1(dp_cluster_1_N171), .A2(n2318), .B(dp_cluster_1_N199), 
        .ZN(n2317) );
  IOA21D1 U2428 ( .A1(n2971), .A2(dp_cluster_3_N116), .B(n2970), .ZN(n2973) );
  OAI21D1 U2429 ( .A1(dp_cluster_3_N116), .A2(n2971), .B(dp_cluster_3_N144), 
        .ZN(n2970) );
  IOA21D1 U2430 ( .A1(n2969), .A2(dp_cluster_3_N115), .B(n2968), .ZN(n2971) );
  OAI21D1 U2431 ( .A1(dp_cluster_3_N115), .A2(n2969), .B(dp_cluster_3_N143), 
        .ZN(n2968) );
  CKBD1 U2432 ( .I(s1_7_r[2]), .Z(n1108) );
  CKBD1 U2433 ( .I(s1_5_r[2]), .Z(n1111) );
  CKBD1 U2434 ( .I(s1_7_i[2]), .Z(n1102) );
  CKBD1 U2435 ( .I(s1_5_i[2]), .Z(n1105) );
  FA1D0 U2436 ( .A(dp_cluster_0_mult_486_C412_n375), .B(
        dp_cluster_0_mult_486_C412_n360), .CI(dp_cluster_0_mult_486_C412_n77), 
        .CO(dp_cluster_0_mult_486_C412_n76), .S(dp_cluster_0_N87) );
  OAI22D1 U2437 ( .A1(n1817), .A2(n1818), .B1(n1816), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n375) );
  NR2D1 U2438 ( .A1(n1802), .A2(n1099), .ZN(dp_cluster_0_mult_486_C412_n360)
         );
  FA1D0 U2439 ( .A(dp_cluster_2_mult_486_C409_n375), .B(
        dp_cluster_2_mult_486_C409_n360), .CI(dp_cluster_2_mult_486_C409_n77), 
        .CO(dp_cluster_2_mult_486_C409_n76), .S(dp_cluster_2_N31) );
  OAI22D1 U2440 ( .A1(n2468), .A2(n2469), .B1(n2467), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n375) );
  NR2D1 U2441 ( .A1(n2453), .A2(n1096), .ZN(dp_cluster_2_mult_486_C409_n360)
         );
  FA1D0 U2442 ( .A(dp_cluster_0_mult_486_C412_n240), .B(
        dp_cluster_0_mult_486_C412_n241), .CI(dp_cluster_0_mult_486_C412_n75), 
        .CO(dp_cluster_0_mult_486_C412_n74), .S(dp_cluster_0_N89) );
  FA1D0 U2443 ( .A(dp_cluster_2_mult_486_C409_n240), .B(
        dp_cluster_2_mult_486_C409_n241), .CI(dp_cluster_2_mult_486_C409_n75), 
        .CO(dp_cluster_2_mult_486_C409_n74), .S(dp_cluster_2_N33) );
  FA1D0 U2444 ( .A(dp_cluster_1_mult_512_C418_n130), .B(
        dp_cluster_1_mult_512_C418_n258), .CI(dp_cluster_1_mult_512_C418_n329), 
        .CO(dp_cluster_1_mult_512_C418_n120), .S(
        dp_cluster_1_mult_512_C418_n121) );
  OAI22D1 U2445 ( .A1(n2179), .A2(n2306), .B1(n2307), .B2(n2178), .ZN(
        dp_cluster_1_mult_512_C418_n258) );
  FA1D0 U2446 ( .A(dp_cluster_1_mult_513_C418_n130), .B(
        dp_cluster_1_mult_513_C418_n258), .CI(dp_cluster_1_mult_513_C418_n329), 
        .CO(dp_cluster_1_mult_513_C418_n120), .S(
        dp_cluster_1_mult_513_C418_n121) );
  OAI22D1 U2447 ( .A1(n2027), .A2(n2154), .B1(n2155), .B2(n2026), .ZN(
        dp_cluster_1_mult_513_C418_n258) );
  FA1D0 U2448 ( .A(dp_cluster_0_mult_486_C412_n130), .B(
        dp_cluster_0_mult_486_C412_n258), .CI(dp_cluster_0_mult_486_C412_n329), 
        .CO(dp_cluster_0_mult_486_C412_n120), .S(
        dp_cluster_0_mult_486_C412_n121) );
  OAI22D1 U2449 ( .A1(n1701), .A2(n1828), .B1(n1829), .B2(n1700), .ZN(
        dp_cluster_0_mult_486_C412_n258) );
  FA1D0 U2450 ( .A(dp_cluster_0_mult_485_C412_n130), .B(
        dp_cluster_0_mult_485_C412_n258), .CI(dp_cluster_0_mult_485_C412_n329), 
        .CO(dp_cluster_0_mult_485_C412_n120), .S(
        dp_cluster_0_mult_485_C412_n121) );
  OAI22D1 U2451 ( .A1(n1853), .A2(n1980), .B1(n1981), .B2(n1852), .ZN(
        dp_cluster_0_mult_485_C412_n258) );
  FA1D0 U2452 ( .A(dp_cluster_3_mult_512_C415_n130), .B(
        dp_cluster_3_mult_512_C415_n258), .CI(dp_cluster_3_mult_512_C415_n329), 
        .CO(dp_cluster_3_mult_512_C415_n120), .S(
        dp_cluster_3_mult_512_C415_n121) );
  OAI22D1 U2453 ( .A1(n2830), .A2(n2957), .B1(n2958), .B2(n2829), .ZN(
        dp_cluster_3_mult_512_C415_n258) );
  FA1D0 U2454 ( .A(dp_cluster_3_mult_513_C415_n130), .B(
        dp_cluster_3_mult_513_C415_n258), .CI(dp_cluster_3_mult_513_C415_n329), 
        .CO(dp_cluster_3_mult_513_C415_n120), .S(
        dp_cluster_3_mult_513_C415_n121) );
  OAI22D1 U2455 ( .A1(n2678), .A2(n2805), .B1(n2806), .B2(n2677), .ZN(
        dp_cluster_3_mult_513_C415_n258) );
  FA1D0 U2456 ( .A(dp_cluster_2_mult_486_C409_n130), .B(
        dp_cluster_2_mult_486_C409_n258), .CI(dp_cluster_2_mult_486_C409_n329), 
        .CO(dp_cluster_2_mult_486_C409_n120), .S(
        dp_cluster_2_mult_486_C409_n121) );
  OAI22D1 U2457 ( .A1(n2352), .A2(n2479), .B1(n2480), .B2(n2351), .ZN(
        dp_cluster_2_mult_486_C409_n258) );
  FA1D0 U2458 ( .A(dp_cluster_2_mult_485_C409_n130), .B(
        dp_cluster_2_mult_485_C409_n258), .CI(dp_cluster_2_mult_485_C409_n329), 
        .CO(dp_cluster_2_mult_485_C409_n120), .S(
        dp_cluster_2_mult_485_C409_n121) );
  OAI22D1 U2459 ( .A1(n2504), .A2(n2631), .B1(n2632), .B2(n2503), .ZN(
        dp_cluster_2_mult_485_C409_n258) );
  XOR3D1 U2460 ( .A1(n1989), .A2(n1988), .A3(n1987), .Z(dp_cluster_0_N84) );
  OAI22D1 U2461 ( .A1(n1986), .A2(n963), .B1(n1984), .B2(n1983), .ZN(n1987) );
  XOR3D1 U2462 ( .A1(n2640), .A2(n2639), .A3(n2638), .Z(dp_cluster_2_N28) );
  OAI22D1 U2463 ( .A1(n2637), .A2(n987), .B1(n2635), .B2(n2634), .ZN(n2638) );
  NR2D1 U2464 ( .A1(dp_cluster_0_N59), .A2(n1993), .ZN(n1992) );
  OAI22D1 U2465 ( .A1(n1991), .A2(n1174), .B1(dp_cluster_0_N86), .B2(n1990), 
        .ZN(n1993) );
  NR2D1 U2466 ( .A1(dp_cluster_2_N3), .A2(n2644), .ZN(n2643) );
  OAI22D1 U2467 ( .A1(n2642), .A2(n1135), .B1(dp_cluster_2_N30), .B2(n2641), 
        .ZN(n2644) );
  CKBD1 U2468 ( .I(n1399), .Z(n1093) );
  CKBD1 U2469 ( .I(n1384), .Z(n1090) );
  CKBD1 U2470 ( .I(s1_7_r[2]), .Z(n1109) );
  CKBD1 U2471 ( .I(s1_5_r[2]), .Z(n1112) );
  CKBD1 U2472 ( .I(s1_7_i[2]), .Z(n1103) );
  CKBD1 U2473 ( .I(s1_5_i[2]), .Z(n1106) );
  INVD1 U2474 ( .I(dp_cluster_0_N60), .ZN(n1171) );
  INVD1 U2475 ( .I(dp_cluster_2_N4), .ZN(n1132) );
  INVD1 U2476 ( .I(dp_cluster_0_N58), .ZN(n1174) );
  INVD1 U2477 ( .I(dp_cluster_2_N2), .ZN(n1135) );
  CKBD1 U2478 ( .I(n1399), .Z(n1094) );
  CKBD1 U2479 ( .I(n1384), .Z(n1091) );
  OAI22D1 U2480 ( .A1(n2280), .A2(n2263), .B1(n2264), .B2(n973), .ZN(
        dp_cluster_1_mult_512_C418_n150) );
  OAI22D1 U2481 ( .A1(n2128), .A2(n2111), .B1(n2112), .B2(n967), .ZN(
        dp_cluster_1_mult_513_C418_n150) );
  OAI22D1 U2482 ( .A1(n1802), .A2(n1785), .B1(n1786), .B2(n955), .ZN(
        dp_cluster_0_mult_486_C412_n150) );
  OAI22D1 U2483 ( .A1(n1954), .A2(n1937), .B1(n1938), .B2(n961), .ZN(
        dp_cluster_0_mult_485_C412_n150) );
  OAI22D1 U2484 ( .A1(n2931), .A2(n2914), .B1(n2915), .B2(n997), .ZN(
        dp_cluster_3_mult_512_C415_n150) );
  OAI22D1 U2485 ( .A1(n2779), .A2(n2762), .B1(n2763), .B2(n991), .ZN(
        dp_cluster_3_mult_513_C415_n150) );
  OAI22D1 U2486 ( .A1(n2453), .A2(n2436), .B1(n2437), .B2(n979), .ZN(
        dp_cluster_2_mult_486_C409_n150) );
  OAI22D1 U2487 ( .A1(n2605), .A2(n2588), .B1(n2589), .B2(n985), .ZN(
        dp_cluster_2_mult_485_C409_n150) );
  OAI22D1 U2488 ( .A1(n2262), .A2(n2245), .B1(n2246), .B2(n972), .ZN(
        dp_cluster_1_mult_512_C418_n130) );
  OAI22D1 U2489 ( .A1(n2110), .A2(n2093), .B1(n2094), .B2(n966), .ZN(
        dp_cluster_1_mult_513_C418_n130) );
  OAI22D1 U2490 ( .A1(n1784), .A2(n1767), .B1(n1768), .B2(n954), .ZN(
        dp_cluster_0_mult_486_C412_n130) );
  OAI22D1 U2491 ( .A1(n1936), .A2(n1919), .B1(n1920), .B2(n960), .ZN(
        dp_cluster_0_mult_485_C412_n130) );
  OAI22D1 U2492 ( .A1(n2913), .A2(n2896), .B1(n2897), .B2(n996), .ZN(
        dp_cluster_3_mult_512_C415_n130) );
  OAI22D1 U2493 ( .A1(n2761), .A2(n2744), .B1(n2745), .B2(n990), .ZN(
        dp_cluster_3_mult_513_C415_n130) );
  OAI22D1 U2494 ( .A1(n2435), .A2(n2418), .B1(n2419), .B2(n978), .ZN(
        dp_cluster_2_mult_486_C409_n130) );
  OAI22D1 U2495 ( .A1(n2587), .A2(n2570), .B1(n2571), .B2(n984), .ZN(
        dp_cluster_2_mult_485_C409_n130) );
  OAI22D1 U2496 ( .A1(n2304), .A2(n2303), .B1(n2302), .B2(n976), .ZN(
        dp_cluster_1_mult_512_C418_n98) );
  OAI22D1 U2497 ( .A1(n2152), .A2(n2151), .B1(n2150), .B2(n970), .ZN(
        dp_cluster_1_mult_513_C418_n98) );
  OAI22D1 U2498 ( .A1(n1826), .A2(n1825), .B1(n1824), .B2(n958), .ZN(
        dp_cluster_0_mult_486_C412_n98) );
  OAI22D1 U2499 ( .A1(n1978), .A2(n1977), .B1(n1976), .B2(n964), .ZN(
        dp_cluster_0_mult_485_C412_n98) );
  OAI22D1 U2500 ( .A1(n2955), .A2(n2954), .B1(n2953), .B2(n1000), .ZN(
        dp_cluster_3_mult_512_C415_n98) );
  OAI22D1 U2501 ( .A1(n2803), .A2(n2802), .B1(n2801), .B2(n994), .ZN(
        dp_cluster_3_mult_513_C415_n98) );
  OAI22D1 U2502 ( .A1(n2477), .A2(n2476), .B1(n2475), .B2(n982), .ZN(
        dp_cluster_2_mult_486_C409_n98) );
  OAI22D1 U2503 ( .A1(n2629), .A2(n2628), .B1(n2627), .B2(n988), .ZN(
        dp_cluster_2_mult_485_C409_n98) );
  OAI22D1 U2504 ( .A1(n2300), .A2(n2299), .B1(n2298), .B2(n971), .ZN(
        dp_cluster_1_mult_512_C418_n86) );
  OAI22D1 U2505 ( .A1(n2148), .A2(n2147), .B1(n2146), .B2(n965), .ZN(
        dp_cluster_1_mult_513_C418_n86) );
  OAI22D1 U2506 ( .A1(n1822), .A2(n1821), .B1(n1820), .B2(n953), .ZN(
        dp_cluster_0_mult_486_C412_n86) );
  OAI22D1 U2507 ( .A1(n1974), .A2(n1973), .B1(n1972), .B2(n959), .ZN(
        dp_cluster_0_mult_485_C412_n86) );
  OAI22D1 U2508 ( .A1(n2951), .A2(n2950), .B1(n2949), .B2(n995), .ZN(
        dp_cluster_3_mult_512_C415_n86) );
  OAI22D1 U2509 ( .A1(n2799), .A2(n2798), .B1(n2797), .B2(n989), .ZN(
        dp_cluster_3_mult_513_C415_n86) );
  OAI22D1 U2510 ( .A1(n2473), .A2(n2472), .B1(n2471), .B2(n977), .ZN(
        dp_cluster_2_mult_486_C409_n86) );
  OAI22D1 U2511 ( .A1(n2625), .A2(n2624), .B1(n2623), .B2(n983), .ZN(
        dp_cluster_2_mult_485_C409_n86) );
  OAI22D1 U2512 ( .A1(n2185), .A2(n975), .B1(n2310), .B2(n2312), .ZN(
        dp_cluster_1_mult_512_C418_n266) );
  OAI22D1 U2513 ( .A1(n2173), .A2(n2306), .B1(n2307), .B2(n2305), .ZN(
        dp_cluster_1_mult_512_C418_n252) );
  OAI22D1 U2514 ( .A1(n2033), .A2(n969), .B1(n2158), .B2(n2160), .ZN(
        dp_cluster_1_mult_513_C418_n266) );
  OAI22D1 U2515 ( .A1(n2021), .A2(n2154), .B1(n2155), .B2(n2153), .ZN(
        dp_cluster_1_mult_513_C418_n252) );
  OAI22D1 U2516 ( .A1(n2836), .A2(n999), .B1(n2961), .B2(n2963), .ZN(
        dp_cluster_3_mult_512_C415_n266) );
  OAI22D1 U2517 ( .A1(n2824), .A2(n2957), .B1(n2958), .B2(n2956), .ZN(
        dp_cluster_3_mult_512_C415_n252) );
  OAI22D1 U2518 ( .A1(n2684), .A2(n993), .B1(n2809), .B2(n2811), .ZN(
        dp_cluster_3_mult_513_C415_n266) );
  OAI22D1 U2519 ( .A1(n2672), .A2(n2805), .B1(n2806), .B2(n2804), .ZN(
        dp_cluster_3_mult_513_C415_n252) );
  OAI22D1 U2520 ( .A1(n1707), .A2(n957), .B1(n1832), .B2(n1834), .ZN(
        dp_cluster_0_mult_486_C412_n266) );
  OAI22D1 U2521 ( .A1(n1695), .A2(n1828), .B1(n1829), .B2(n1827), .ZN(
        dp_cluster_0_mult_486_C412_n252) );
  OAI22D1 U2522 ( .A1(n1859), .A2(n963), .B1(n1984), .B2(n1986), .ZN(
        dp_cluster_0_mult_485_C412_n266) );
  OAI22D1 U2523 ( .A1(n1847), .A2(n1980), .B1(n1981), .B2(n1979), .ZN(
        dp_cluster_0_mult_485_C412_n252) );
  OAI22D1 U2524 ( .A1(n2358), .A2(n981), .B1(n2483), .B2(n2485), .ZN(
        dp_cluster_2_mult_486_C409_n266) );
  OAI22D1 U2525 ( .A1(n2346), .A2(n2479), .B1(n2480), .B2(n2478), .ZN(
        dp_cluster_2_mult_486_C409_n252) );
  OAI22D1 U2526 ( .A1(n2510), .A2(n987), .B1(n2635), .B2(n2637), .ZN(
        dp_cluster_2_mult_485_C409_n266) );
  OAI22D1 U2527 ( .A1(n2498), .A2(n2631), .B1(n2632), .B2(n2630), .ZN(
        dp_cluster_2_mult_485_C409_n252) );
  ND2D1 U2528 ( .A1(s2_5_i[0]), .A2(n939), .ZN(sub_383_carry[1]) );
  INVD1 U2529 ( .I(s2_5_i[1]), .ZN(n1634) );
  INVD1 U2530 ( .I(s2_4_i[0]), .ZN(n939) );
  INVD1 U2531 ( .I(s2_5_i[2]), .ZN(n1632) );
  INVD1 U2532 ( .I(s2_5_i[3]), .ZN(n1630) );
  INVD1 U2533 ( .I(s2_5_i[4]), .ZN(n1628) );
  INVD1 U2534 ( .I(s2_5_i[5]), .ZN(n1626) );
  INVD1 U2535 ( .I(s2_5_i[6]), .ZN(n1624) );
  INVD1 U2536 ( .I(s2_5_i[7]), .ZN(n1622) );
  INVD1 U2537 ( .I(s2_5_i[8]), .ZN(n1620) );
  INVD1 U2538 ( .I(s2_5_i[9]), .ZN(n1618) );
  INVD1 U2539 ( .I(s2_5_i[10]), .ZN(n1616) );
  INVD1 U2540 ( .I(s2_5_i[11]), .ZN(n1614) );
  INVD1 U2541 ( .I(s2_5_i[12]), .ZN(n1612) );
  INVD1 U2542 ( .I(s2_5_i[13]), .ZN(n1610) );
  INVD1 U2543 ( .I(s2_5_i[14]), .ZN(n1608) );
  ND2D1 U2544 ( .A1(s2_5_r[0]), .A2(n943), .ZN(sub_374_carry[1]) );
  INVD1 U2545 ( .I(s2_5_r[1]), .ZN(n1600) );
  INVD1 U2546 ( .I(s2_4_r[0]), .ZN(n943) );
  INVD1 U2547 ( .I(s2_5_r[2]), .ZN(n1597) );
  INVD1 U2548 ( .I(s2_5_r[3]), .ZN(n1594) );
  INVD1 U2549 ( .I(s2_5_r[4]), .ZN(n1591) );
  INVD1 U2550 ( .I(s2_5_r[5]), .ZN(n1588) );
  INVD1 U2551 ( .I(s2_5_r[6]), .ZN(n1585) );
  INVD1 U2552 ( .I(s2_5_r[7]), .ZN(n1582) );
  INVD1 U2553 ( .I(s2_5_r[8]), .ZN(n1579) );
  INVD1 U2554 ( .I(s2_5_r[9]), .ZN(n1576) );
  INVD1 U2555 ( .I(s2_5_r[10]), .ZN(n1573) );
  INVD1 U2556 ( .I(s2_5_r[11]), .ZN(n1570) );
  INVD1 U2557 ( .I(s2_5_r[12]), .ZN(n1567) );
  INVD1 U2558 ( .I(s2_5_r[13]), .ZN(n1564) );
  INVD1 U2559 ( .I(s2_5_r[14]), .ZN(n1561) );
  ND2D1 U2560 ( .A1(s2_3_tmp_i_0_), .A2(n940), .ZN(sub_381_carry[1]) );
  INVD1 U2561 ( .I(dp_cluster_5_s2_3_r[9]), .ZN(n1473) );
  INVD1 U2562 ( .I(s2_2_i[0]), .ZN(n940) );
  INVD1 U2563 ( .I(dp_cluster_5_s2_3_r[2]), .ZN(n1452) );
  INVD1 U2564 ( .I(dp_cluster_5_s2_3_r[1]), .ZN(n1449) );
  INVD1 U2565 ( .I(dp_cluster_5_s2_3_r[15]), .ZN(n1446) );
  INVD1 U2566 ( .I(dp_cluster_5_s2_3_r[14]), .ZN(n1443) );
  INVD1 U2567 ( .I(dp_cluster_5_s2_3_r[13]), .ZN(n1440) );
  INVD1 U2568 ( .I(dp_cluster_5_s2_3_r[12]), .ZN(n1437) );
  INVD1 U2569 ( .I(dp_cluster_5_s2_3_r[11]), .ZN(n1434) );
  ND2D1 U2570 ( .A1(s2_3_i[0]), .A2(n944), .ZN(sub_372_carry[1]) );
  INVD1 U2571 ( .I(s2_3_i[1]), .ZN(n1507) );
  INVD1 U2572 ( .I(s2_2_r[0]), .ZN(n944) );
  INVD1 U2573 ( .I(s2_3_i[2]), .ZN(n1505) );
  INVD1 U2574 ( .I(s2_3_i[3]), .ZN(n1503) );
  INVD1 U2575 ( .I(s2_3_i[4]), .ZN(n1501) );
  INVD1 U2576 ( .I(s2_3_i[5]), .ZN(n1499) );
  INVD1 U2577 ( .I(s2_3_i[6]), .ZN(n1497) );
  INVD1 U2578 ( .I(s2_3_i[7]), .ZN(n1495) );
  INVD1 U2579 ( .I(s2_3_i[8]), .ZN(n1493) );
  INVD1 U2580 ( .I(s2_3_i[9]), .ZN(n1491) );
  INVD1 U2581 ( .I(s2_3_i[10]), .ZN(n1489) );
  INVD1 U2582 ( .I(s2_3_i[11]), .ZN(n1487) );
  INVD1 U2583 ( .I(s2_3_i[12]), .ZN(n1485) );
  INVD1 U2584 ( .I(s2_3_i[13]), .ZN(n1483) );
  INVD1 U2585 ( .I(s2_3_i[14]), .ZN(n1481) );
  ND2D1 U2586 ( .A1(s2_1_i[0]), .A2(n941), .ZN(sub_379_carry[1]) );
  INVD1 U2587 ( .I(s2_1_i[1]), .ZN(n1506) );
  INVD1 U2588 ( .I(s2_0_i[0]), .ZN(n941) );
  INVD1 U2589 ( .I(s2_1_i[2]), .ZN(n1504) );
  INVD1 U2590 ( .I(s2_1_i[3]), .ZN(n1502) );
  INVD1 U2591 ( .I(s2_1_i[4]), .ZN(n1500) );
  INVD1 U2592 ( .I(s2_1_i[5]), .ZN(n1498) );
  INVD1 U2593 ( .I(s2_1_i[6]), .ZN(n1496) );
  INVD1 U2594 ( .I(s2_1_i[7]), .ZN(n1494) );
  INVD1 U2595 ( .I(s2_1_i[8]), .ZN(n1492) );
  INVD1 U2596 ( .I(s2_1_i[9]), .ZN(n1490) );
  INVD1 U2597 ( .I(s2_1_i[10]), .ZN(n1488) );
  INVD1 U2598 ( .I(s2_1_i[11]), .ZN(n1486) );
  INVD1 U2599 ( .I(s2_1_i[12]), .ZN(n1484) );
  INVD1 U2600 ( .I(s2_1_i[13]), .ZN(n1482) );
  INVD1 U2601 ( .I(s2_1_i[14]), .ZN(n1480) );
  ND2D1 U2602 ( .A1(s2_1_r[0]), .A2(n945), .ZN(sub_370_carry[1]) );
  INVD1 U2603 ( .I(s2_1_r[1]), .ZN(n1472) );
  INVD1 U2604 ( .I(s2_0_r[0]), .ZN(n945) );
  INVD1 U2605 ( .I(s2_1_r[2]), .ZN(n1469) );
  INVD1 U2606 ( .I(s2_1_r[3]), .ZN(n1466) );
  INVD1 U2607 ( .I(s2_1_r[4]), .ZN(n1463) );
  INVD1 U2608 ( .I(s2_1_r[5]), .ZN(n1460) );
  INVD1 U2609 ( .I(s2_1_r[6]), .ZN(n1457) );
  INVD1 U2610 ( .I(s2_1_r[7]), .ZN(n1454) );
  INVD1 U2611 ( .I(s2_1_r[8]), .ZN(n1451) );
  INVD1 U2612 ( .I(s2_1_r[9]), .ZN(n1448) );
  INVD1 U2613 ( .I(s2_1_r[10]), .ZN(n1445) );
  INVD1 U2614 ( .I(s2_1_r[11]), .ZN(n1442) );
  INVD1 U2615 ( .I(s2_1_r[12]), .ZN(n1439) );
  INVD1 U2616 ( .I(s2_1_r[13]), .ZN(n1436) );
  INVD1 U2617 ( .I(s2_1_r[14]), .ZN(n1433) );
  INVD1 U2618 ( .I(s2_7_i[14]), .ZN(n1609) );
  INVD1 U2619 ( .I(s2_7_i[13]), .ZN(n1611) );
  INVD1 U2620 ( .I(s2_7_i[12]), .ZN(n1613) );
  INVD1 U2621 ( .I(s2_7_i[11]), .ZN(n1615) );
  INVD1 U2622 ( .I(s2_7_i[10]), .ZN(n1617) );
  INVD1 U2623 ( .I(s2_7_i[9]), .ZN(n1619) );
  INVD1 U2624 ( .I(s2_7_i[8]), .ZN(n1621) );
  INVD1 U2625 ( .I(s2_7_i[7]), .ZN(n1623) );
  INVD1 U2626 ( .I(s2_7_i[6]), .ZN(n1625) );
  INVD1 U2627 ( .I(s2_7_i[5]), .ZN(n1627) );
  INVD1 U2628 ( .I(s2_7_i[4]), .ZN(n1629) );
  INVD1 U2629 ( .I(s2_7_i[3]), .ZN(n1631) );
  INVD1 U2630 ( .I(s2_7_i[2]), .ZN(n1633) );
  ND2D1 U2631 ( .A1(s2_7_i[0]), .A2(n942), .ZN(sub_376_carry[1]) );
  INVD1 U2632 ( .I(s2_7_i[1]), .ZN(n1635) );
  INVD1 U2633 ( .I(s2_6_r[0]), .ZN(n942) );
  INVD1 U2634 ( .I(dp_cluster_4_s2_7_r[11]), .ZN(n1562) );
  INVD1 U2635 ( .I(dp_cluster_4_s2_7_r[12]), .ZN(n1565) );
  INVD1 U2636 ( .I(dp_cluster_4_s2_7_r[13]), .ZN(n1568) );
  INVD1 U2637 ( .I(dp_cluster_4_s2_7_r[14]), .ZN(n1571) );
  INVD1 U2638 ( .I(dp_cluster_4_s2_7_r[15]), .ZN(n1574) );
  INVD1 U2639 ( .I(dp_cluster_4_s2_7_r[1]), .ZN(n1577) );
  INVD1 U2640 ( .I(dp_cluster_4_s2_7_r[2]), .ZN(n1580) );
  ND2D1 U2641 ( .A1(s2_7_tmp_i_0_), .A2(n938), .ZN(sub_385_carry[1]) );
  INVD1 U2642 ( .I(dp_cluster_4_s2_7_r[9]), .ZN(n1601) );
  INVD1 U2643 ( .I(s2_6_i[0]), .ZN(n938) );
  FA1D0 U2644 ( .A(dp_cluster_1_mult_512_C418_n268), .B(
        dp_cluster_1_mult_512_C418_n254), .CI(dp_cluster_1_mult_512_C418_n296), 
        .CO(dp_cluster_1_mult_512_C418_n91), .S(dp_cluster_1_mult_512_C418_n92) );
  OAI22D1 U2645 ( .A1(n2187), .A2(n975), .B1(n2310), .B2(n2186), .ZN(
        dp_cluster_1_mult_512_C418_n268) );
  OAI22D1 U2646 ( .A1(n2175), .A2(n2306), .B1(n2307), .B2(n2174), .ZN(
        dp_cluster_1_mult_512_C418_n254) );
  FA1D0 U2647 ( .A(dp_cluster_1_mult_513_C418_n268), .B(
        dp_cluster_1_mult_513_C418_n254), .CI(dp_cluster_1_mult_513_C418_n296), 
        .CO(dp_cluster_1_mult_513_C418_n91), .S(dp_cluster_1_mult_513_C418_n92) );
  OAI22D1 U2648 ( .A1(n2035), .A2(n969), .B1(n2158), .B2(n2034), .ZN(
        dp_cluster_1_mult_513_C418_n268) );
  OAI22D1 U2649 ( .A1(n2023), .A2(n2154), .B1(n2155), .B2(n2022), .ZN(
        dp_cluster_1_mult_513_C418_n254) );
  FA1D0 U2650 ( .A(dp_cluster_0_mult_486_C412_n268), .B(
        dp_cluster_0_mult_486_C412_n254), .CI(dp_cluster_0_mult_486_C412_n296), 
        .CO(dp_cluster_0_mult_486_C412_n91), .S(dp_cluster_0_mult_486_C412_n92) );
  OAI22D1 U2651 ( .A1(n1709), .A2(n957), .B1(n1832), .B2(n1708), .ZN(
        dp_cluster_0_mult_486_C412_n268) );
  OAI22D1 U2652 ( .A1(n1697), .A2(n1828), .B1(n1829), .B2(n1696), .ZN(
        dp_cluster_0_mult_486_C412_n254) );
  FA1D0 U2653 ( .A(dp_cluster_0_mult_485_C412_n268), .B(
        dp_cluster_0_mult_485_C412_n254), .CI(dp_cluster_0_mult_485_C412_n296), 
        .CO(dp_cluster_0_mult_485_C412_n91), .S(dp_cluster_0_mult_485_C412_n92) );
  OAI22D1 U2654 ( .A1(n1861), .A2(n963), .B1(n1984), .B2(n1860), .ZN(
        dp_cluster_0_mult_485_C412_n268) );
  OAI22D1 U2655 ( .A1(n1849), .A2(n1980), .B1(n1981), .B2(n1848), .ZN(
        dp_cluster_0_mult_485_C412_n254) );
  FA1D0 U2656 ( .A(dp_cluster_3_mult_512_C415_n268), .B(
        dp_cluster_3_mult_512_C415_n254), .CI(dp_cluster_3_mult_512_C415_n296), 
        .CO(dp_cluster_3_mult_512_C415_n91), .S(dp_cluster_3_mult_512_C415_n92) );
  OAI22D1 U2657 ( .A1(n2838), .A2(n999), .B1(n2961), .B2(n2837), .ZN(
        dp_cluster_3_mult_512_C415_n268) );
  OAI22D1 U2658 ( .A1(n2826), .A2(n2957), .B1(n2958), .B2(n2825), .ZN(
        dp_cluster_3_mult_512_C415_n254) );
  FA1D0 U2659 ( .A(dp_cluster_3_mult_513_C415_n268), .B(
        dp_cluster_3_mult_513_C415_n254), .CI(dp_cluster_3_mult_513_C415_n296), 
        .CO(dp_cluster_3_mult_513_C415_n91), .S(dp_cluster_3_mult_513_C415_n92) );
  OAI22D1 U2660 ( .A1(n2686), .A2(n993), .B1(n2809), .B2(n2685), .ZN(
        dp_cluster_3_mult_513_C415_n268) );
  OAI22D1 U2661 ( .A1(n2674), .A2(n2805), .B1(n2806), .B2(n2673), .ZN(
        dp_cluster_3_mult_513_C415_n254) );
  FA1D0 U2662 ( .A(dp_cluster_2_mult_486_C409_n268), .B(
        dp_cluster_2_mult_486_C409_n254), .CI(dp_cluster_2_mult_486_C409_n296), 
        .CO(dp_cluster_2_mult_486_C409_n91), .S(dp_cluster_2_mult_486_C409_n92) );
  OAI22D1 U2663 ( .A1(n2360), .A2(n981), .B1(n2483), .B2(n2359), .ZN(
        dp_cluster_2_mult_486_C409_n268) );
  OAI22D1 U2664 ( .A1(n2348), .A2(n2479), .B1(n2480), .B2(n2347), .ZN(
        dp_cluster_2_mult_486_C409_n254) );
  FA1D0 U2665 ( .A(dp_cluster_2_mult_485_C409_n268), .B(
        dp_cluster_2_mult_485_C409_n254), .CI(dp_cluster_2_mult_485_C409_n296), 
        .CO(dp_cluster_2_mult_485_C409_n91), .S(dp_cluster_2_mult_485_C409_n92) );
  OAI22D1 U2666 ( .A1(n2512), .A2(n987), .B1(n2635), .B2(n2511), .ZN(
        dp_cluster_2_mult_485_C409_n268) );
  OAI22D1 U2667 ( .A1(n2500), .A2(n2631), .B1(n2632), .B2(n2499), .ZN(
        dp_cluster_2_mult_485_C409_n254) );
  IOA21D1 U2668 ( .A1(dp_cluster_1_N170), .A2(dp_cluster_1_N198), .B(n2316), 
        .ZN(n2318) );
  OAI211D1 U2669 ( .A1(dp_cluster_1_N170), .A2(dp_cluster_1_N198), .B(
        dp_cluster_1_N169), .C(dp_cluster_1_N197), .ZN(n2316) );
  NR2D1 U2670 ( .A1(n1044), .A2(n1099), .ZN(dp_cluster_1_N169) );
  NR2D1 U2671 ( .A1(n1088), .A2(n1093), .ZN(dp_cluster_1_N197) );
  IOA21D1 U2672 ( .A1(dp_cluster_3_N114), .A2(dp_cluster_3_N142), .B(n2967), 
        .ZN(n2969) );
  OAI211D1 U2673 ( .A1(dp_cluster_3_N114), .A2(dp_cluster_3_N142), .B(
        dp_cluster_3_N113), .C(dp_cluster_3_N141), .ZN(n2967) );
  NR2D1 U2674 ( .A1(n1022), .A2(n1096), .ZN(dp_cluster_3_N113) );
  NR2D1 U2675 ( .A1(n1066), .A2(n1090), .ZN(dp_cluster_3_N141) );
  CKXOR2D1 U2676 ( .A1(s1_6_r[16]), .A2(n952), .Z(s1_6_tmp_i[15]) );
  ND2D1 U2677 ( .A1(n933), .A2(n1137), .ZN(n952) );
  INVD1 U2678 ( .I(s2_5_i[0]), .ZN(n1636) );
  INVD1 U2679 ( .I(s2_5_r[0]), .ZN(n1603) );
  INVD1 U2680 ( .I(s2_1_i[0]), .ZN(n1508) );
  INVD1 U2681 ( .I(s2_1_r[0]), .ZN(n1475) );
  INVD1 U2682 ( .I(s2_3_i[0]), .ZN(n1509) );
  INVD1 U2683 ( .I(s2_7_i[0]), .ZN(n1637) );
  INVD1 U2684 ( .I(s2_3_tmp_i_0_), .ZN(n1476) );
  INVD1 U2685 ( .I(s2_7_tmp_i_0_), .ZN(n1604) );
  INVD1 U2686 ( .I(s2_5_i[15]), .ZN(n1606) );
  INVD1 U2687 ( .I(s2_5_r[15]), .ZN(n1558) );
  INVD1 U2688 ( .I(dp_cluster_5_s2_3_r[10]), .ZN(n1431) );
  INVD1 U2689 ( .I(s2_3_i[15]), .ZN(n1479) );
  INVD1 U2690 ( .I(s2_1_i[15]), .ZN(n1478) );
  INVD1 U2691 ( .I(s2_1_r[15]), .ZN(n1430) );
  INVD1 U2692 ( .I(s2_7_i[15]), .ZN(n1607) );
  INVD1 U2693 ( .I(dp_cluster_4_s2_7_r[10]), .ZN(n1559) );
  CKBD1 U2694 ( .I(n1399), .Z(n1092) );
  CKBD1 U2695 ( .I(n1384), .Z(n1089) );
  CKBD1 U2696 ( .I(n1429), .Z(n1098) );
  CKBD1 U2697 ( .I(n1414), .Z(n1095) );
  CKBD1 U2698 ( .I(n1429), .Z(n1099) );
  CKBD1 U2699 ( .I(n1414), .Z(n1096) );
  INVD1 U2700 ( .I(s1_6_r[4]), .ZN(n1148) );
  INVD1 U2701 ( .I(s1_6_r[5]), .ZN(n1147) );
  INVD1 U2702 ( .I(s1_6_r[6]), .ZN(n1146) );
  INVD1 U2703 ( .I(s1_6_r[7]), .ZN(n1145) );
  INVD1 U2704 ( .I(s1_6_r[8]), .ZN(n1144) );
  INVD1 U2705 ( .I(s1_6_r[9]), .ZN(n1143) );
  INVD1 U2706 ( .I(s1_6_r[10]), .ZN(n1142) );
  INVD1 U2707 ( .I(s1_6_r[11]), .ZN(n1141) );
  INVD1 U2708 ( .I(s1_6_r[12]), .ZN(n1140) );
  INVD1 U2709 ( .I(s1_6_r[13]), .ZN(n1139) );
  INVD1 U2710 ( .I(s1_6_r[14]), .ZN(n1138) );
  INVD1 U2711 ( .I(s1_6_r[15]), .ZN(n1137) );
  CKBD1 U2712 ( .I(n1429), .Z(n1100) );
  CKBD1 U2713 ( .I(n1414), .Z(n1097) );
  INVD1 U2714 ( .I(dp_cluster_5_s2_3_r[8]), .ZN(n1470) );
  INVD1 U2715 ( .I(dp_cluster_5_s2_3_r[7]), .ZN(n1467) );
  INVD1 U2716 ( .I(dp_cluster_5_s2_3_r[6]), .ZN(n1464) );
  INVD1 U2717 ( .I(dp_cluster_5_s2_3_r[5]), .ZN(n1461) );
  INVD1 U2718 ( .I(dp_cluster_5_s2_3_r[4]), .ZN(n1458) );
  INVD1 U2719 ( .I(dp_cluster_5_s2_3_r[3]), .ZN(n1455) );
  INVD1 U2720 ( .I(dp_cluster_4_s2_7_r[3]), .ZN(n1583) );
  INVD1 U2721 ( .I(dp_cluster_4_s2_7_r[4]), .ZN(n1586) );
  INVD1 U2722 ( .I(dp_cluster_4_s2_7_r[5]), .ZN(n1589) );
  INVD1 U2723 ( .I(dp_cluster_4_s2_7_r[6]), .ZN(n1592) );
  INVD1 U2724 ( .I(dp_cluster_4_s2_7_r[7]), .ZN(n1595) );
  INVD1 U2725 ( .I(dp_cluster_4_s2_7_r[8]), .ZN(n1598) );
  INVD1 U2726 ( .I(s1_6_tmp_i[0]), .ZN(n1151) );
  INVD1 U2727 ( .I(s1_6_r[2]), .ZN(n1150) );
  INVD1 U2728 ( .I(s1_6_r[3]), .ZN(n1149) );
  HA1D0 U2729 ( .A(dp_cluster_0_mult_485_C412_n247), .B(
        dp_cluster_0_mult_485_C412_n327), .CO(dp_cluster_0_mult_485_C412_n230), 
        .S(dp_cluster_0_mult_485_C412_n231) );
  OAI22D1 U2730 ( .A1(n1917), .A2(n962), .B1(n1918), .B2(n1915), .ZN(
        dp_cluster_0_mult_485_C412_n327) );
  OAI32D1 U2731 ( .A1(n1033), .A2(W3_8_r[48]), .A3(n1918), .B1(n1033), .B2(
        n962), .ZN(dp_cluster_0_mult_485_C412_n247) );
  HA1D0 U2732 ( .A(dp_cluster_2_mult_485_C409_n247), .B(
        dp_cluster_2_mult_485_C409_n327), .CO(dp_cluster_2_mult_485_C409_n230), 
        .S(dp_cluster_2_mult_485_C409_n231) );
  OAI22D1 U2733 ( .A1(n2568), .A2(n986), .B1(n2569), .B2(n2566), .ZN(
        dp_cluster_2_mult_485_C409_n327) );
  OAI32D1 U2734 ( .A1(n1011), .A2(W1_8_r[48]), .A3(n2569), .B1(n1011), .B2(
        n986), .ZN(dp_cluster_2_mult_485_C409_n247) );
  HA1D0 U2735 ( .A(dp_cluster_0_mult_486_C412_n247), .B(
        dp_cluster_0_mult_486_C412_n327), .CO(dp_cluster_0_mult_486_C412_n230), 
        .S(dp_cluster_0_mult_486_C412_n231) );
  OAI22D1 U2736 ( .A1(n1765), .A2(n956), .B1(n1766), .B2(n1763), .ZN(
        dp_cluster_0_mult_486_C412_n327) );
  OAI32D1 U2737 ( .A1(n1077), .A2(W3_8_i[48]), .A3(n1766), .B1(n1077), .B2(
        n956), .ZN(dp_cluster_0_mult_486_C412_n247) );
  HA1D0 U2738 ( .A(dp_cluster_2_mult_486_C409_n247), .B(
        dp_cluster_2_mult_486_C409_n327), .CO(dp_cluster_2_mult_486_C409_n230), 
        .S(dp_cluster_2_mult_486_C409_n231) );
  OAI22D1 U2739 ( .A1(n2416), .A2(n980), .B1(n2417), .B2(n2414), .ZN(
        dp_cluster_2_mult_486_C409_n327) );
  OAI32D1 U2740 ( .A1(n1055), .A2(W1_8_i[48]), .A3(n2417), .B1(n1055), .B2(
        n980), .ZN(dp_cluster_2_mult_486_C409_n247) );
  HA1D0 U2741 ( .A(dp_cluster_1_mult_512_C418_n243), .B(
        dp_cluster_1_mult_512_C418_n263), .CO(dp_cluster_1_mult_512_C418_n172), 
        .S(dp_cluster_1_mult_512_C418_n173) );
  OAI22D1 U2742 ( .A1(n2184), .A2(n2306), .B1(n2307), .B2(n2183), .ZN(
        dp_cluster_1_mult_512_C418_n263) );
  OAI32D1 U2743 ( .A1(n1023), .A2(W3_8_i[48]), .A3(n2307), .B1(n1023), .B2(
        n2306), .ZN(dp_cluster_1_mult_512_C418_n243) );
  HA1D0 U2744 ( .A(dp_cluster_1_mult_513_C418_n243), .B(
        dp_cluster_1_mult_513_C418_n263), .CO(dp_cluster_1_mult_513_C418_n172), 
        .S(dp_cluster_1_mult_513_C418_n173) );
  OAI22D1 U2745 ( .A1(n2032), .A2(n2154), .B1(n2155), .B2(n2031), .ZN(
        dp_cluster_1_mult_513_C418_n263) );
  OAI32D1 U2746 ( .A1(n1067), .A2(W3_8_r[48]), .A3(n2155), .B1(n1067), .B2(
        n2154), .ZN(dp_cluster_1_mult_513_C418_n243) );
  HA1D0 U2747 ( .A(dp_cluster_3_mult_512_C415_n243), .B(
        dp_cluster_3_mult_512_C415_n263), .CO(dp_cluster_3_mult_512_C415_n172), 
        .S(dp_cluster_3_mult_512_C415_n173) );
  OAI22D1 U2748 ( .A1(n2835), .A2(n2957), .B1(n2958), .B2(n2834), .ZN(
        dp_cluster_3_mult_512_C415_n263) );
  OAI32D1 U2749 ( .A1(n1001), .A2(W1_8_i[48]), .A3(n2958), .B1(n1001), .B2(
        n2957), .ZN(dp_cluster_3_mult_512_C415_n243) );
  HA1D0 U2750 ( .A(dp_cluster_3_mult_513_C415_n243), .B(
        dp_cluster_3_mult_513_C415_n263), .CO(dp_cluster_3_mult_513_C415_n172), 
        .S(dp_cluster_3_mult_513_C415_n173) );
  OAI22D1 U2751 ( .A1(n2683), .A2(n2805), .B1(n2806), .B2(n2682), .ZN(
        dp_cluster_3_mult_513_C415_n263) );
  OAI32D1 U2752 ( .A1(n1045), .A2(W1_8_r[48]), .A3(n2806), .B1(n1045), .B2(
        n2805), .ZN(dp_cluster_3_mult_513_C415_n243) );
  INVD1 U2753 ( .I(xi7_i[63]), .ZN(n1354) );
  INVD1 U2754 ( .I(xi5_i[63]), .ZN(n1322) );
  INVD1 U2755 ( .I(xi7_r[63]), .ZN(n1224) );
  INVD1 U2756 ( .I(xi5_r[63]), .ZN(n1192) );
  HA1D0 U2757 ( .A(dp_cluster_1_mult_512_C418_n376), .B(
        dp_cluster_1_mult_512_C418_n250), .CO(dp_cluster_1_mult_512_C418_n77), 
        .S(dp_cluster_1_N170) );
  IOA21D1 U2758 ( .A1(n1100), .A2(n1109), .B(n2296), .ZN(
        dp_cluster_1_mult_512_C418_n250) );
  OAI22D1 U2759 ( .A1(W3_8_i[48]), .A2(n2296), .B1(n2295), .B2(n1042), .ZN(
        dp_cluster_1_mult_512_C418_n376) );
  HA1D0 U2760 ( .A(dp_cluster_1_mult_513_C418_n376), .B(
        dp_cluster_1_mult_513_C418_n250), .CO(dp_cluster_1_mult_513_C418_n77), 
        .S(dp_cluster_1_N198) );
  IOA21D1 U2761 ( .A1(n1094), .A2(n1103), .B(n2144), .ZN(
        dp_cluster_1_mult_513_C418_n250) );
  OAI22D1 U2762 ( .A1(W3_8_r[48]), .A2(n2144), .B1(n2143), .B2(n1086), .ZN(
        dp_cluster_1_mult_513_C418_n376) );
  HA1D0 U2763 ( .A(dp_cluster_3_mult_512_C415_n376), .B(
        dp_cluster_3_mult_512_C415_n250), .CO(dp_cluster_3_mult_512_C415_n77), 
        .S(dp_cluster_3_N114) );
  IOA21D1 U2764 ( .A1(n1097), .A2(n1112), .B(n2947), .ZN(
        dp_cluster_3_mult_512_C415_n250) );
  OAI22D1 U2765 ( .A1(W1_8_i[48]), .A2(n2947), .B1(n2946), .B2(n1020), .ZN(
        dp_cluster_3_mult_512_C415_n376) );
  HA1D0 U2766 ( .A(dp_cluster_3_mult_513_C415_n376), .B(
        dp_cluster_3_mult_513_C415_n250), .CO(dp_cluster_3_mult_513_C415_n77), 
        .S(dp_cluster_3_N142) );
  IOA21D1 U2767 ( .A1(n1091), .A2(n1106), .B(n2795), .ZN(
        dp_cluster_3_mult_513_C415_n250) );
  OAI22D1 U2768 ( .A1(W1_8_r[48]), .A2(n2795), .B1(n2794), .B2(n1064), .ZN(
        dp_cluster_3_mult_513_C415_n376) );
  HA1D0 U2769 ( .A(dp_cluster_0_mult_486_C412_n376), .B(
        dp_cluster_0_mult_486_C412_n250), .CO(dp_cluster_0_mult_486_C412_n77), 
        .S(dp_cluster_0_N86) );
  IOA21D1 U2770 ( .A1(n1100), .A2(n1103), .B(n1818), .ZN(
        dp_cluster_0_mult_486_C412_n250) );
  OAI22D1 U2771 ( .A1(W3_8_i[48]), .A2(n1818), .B1(n1817), .B2(n1087), .ZN(
        dp_cluster_0_mult_486_C412_n376) );
  HA1D0 U2772 ( .A(dp_cluster_2_mult_486_C409_n376), .B(
        dp_cluster_2_mult_486_C409_n250), .CO(dp_cluster_2_mult_486_C409_n77), 
        .S(dp_cluster_2_N30) );
  IOA21D1 U2773 ( .A1(n1097), .A2(n1106), .B(n2469), .ZN(
        dp_cluster_2_mult_486_C409_n250) );
  OAI22D1 U2774 ( .A1(W1_8_i[48]), .A2(n2469), .B1(n2468), .B2(n1065), .ZN(
        dp_cluster_2_mult_486_C409_n376) );
  INVD1 U2775 ( .I(W3_8_r[48]), .ZN(n1399) );
  INVD1 U2776 ( .I(W1_8_r[48]), .ZN(n1384) );
  FA1D0 U2777 ( .A(dp_cluster_1_mult_513_C418_n242), .B(
        dp_cluster_1_mult_513_C418_n249), .CI(dp_cluster_1_mult_513_C418_n76), 
        .CO(dp_cluster_1_mult_513_C418_n75), .S(dp_cluster_1_N200) );
  OAI32D1 U2778 ( .A1(n1083), .A2(W3_8_r[48]), .A3(n2128), .B1(n1083), .B2(
        n967), .ZN(dp_cluster_1_mult_513_C418_n249) );
  FA1D0 U2779 ( .A(dp_cluster_3_mult_513_C415_n242), .B(
        dp_cluster_3_mult_513_C415_n249), .CI(dp_cluster_3_mult_513_C415_n76), 
        .CO(dp_cluster_3_mult_513_C415_n75), .S(dp_cluster_3_N144) );
  OAI32D1 U2780 ( .A1(n1061), .A2(W1_8_r[48]), .A3(n2779), .B1(n1061), .B2(
        n991), .ZN(dp_cluster_3_mult_513_C415_n249) );
  FA1D0 U2781 ( .A(dp_cluster_1_mult_512_C418_n242), .B(
        dp_cluster_1_mult_512_C418_n249), .CI(dp_cluster_1_mult_512_C418_n76), 
        .CO(dp_cluster_1_mult_512_C418_n75), .S(dp_cluster_1_N172) );
  OAI32D1 U2782 ( .A1(n1039), .A2(W3_8_i[48]), .A3(n2280), .B1(n1039), .B2(
        n973), .ZN(dp_cluster_1_mult_512_C418_n249) );
  FA1D0 U2783 ( .A(dp_cluster_3_mult_512_C415_n242), .B(
        dp_cluster_3_mult_512_C415_n249), .CI(dp_cluster_3_mult_512_C415_n76), 
        .CO(dp_cluster_3_mult_512_C415_n75), .S(dp_cluster_3_N116) );
  OAI32D1 U2784 ( .A1(n1017), .A2(W1_8_i[48]), .A3(n2931), .B1(n1017), .B2(
        n997), .ZN(dp_cluster_3_mult_512_C415_n249) );
  FA1D0 U2785 ( .A(dp_cluster_0_mult_486_C412_n242), .B(
        dp_cluster_0_mult_486_C412_n249), .CI(dp_cluster_0_mult_486_C412_n76), 
        .CO(dp_cluster_0_mult_486_C412_n75), .S(dp_cluster_0_N88) );
  OAI32D1 U2786 ( .A1(n1083), .A2(W3_8_i[48]), .A3(n1802), .B1(n1083), .B2(
        n955), .ZN(dp_cluster_0_mult_486_C412_n249) );
  FA1D0 U2787 ( .A(dp_cluster_2_mult_486_C409_n242), .B(
        dp_cluster_2_mult_486_C409_n249), .CI(dp_cluster_2_mult_486_C409_n76), 
        .CO(dp_cluster_2_mult_486_C409_n75), .S(dp_cluster_2_N32) );
  OAI32D1 U2788 ( .A1(n1061), .A2(W1_8_i[48]), .A3(n2453), .B1(n1061), .B2(
        n979), .ZN(dp_cluster_2_mult_486_C409_n249) );
  INVD1 U2789 ( .I(xi7_r[49]), .ZN(n1238) );
  INVD1 U2790 ( .I(xi5_r[49]), .ZN(n1206) );
  INVD1 U2791 ( .I(xi7_i[49]), .ZN(n1368) );
  INVD1 U2792 ( .I(xi5_i[49]), .ZN(n1336) );
  INVD1 U2793 ( .I(xi7_i[50]), .ZN(n1367) );
  INVD1 U2794 ( .I(xi7_r[50]), .ZN(n1237) );
  INVD1 U2795 ( .I(xi5_i[50]), .ZN(n1335) );
  INVD1 U2796 ( .I(xi5_r[50]), .ZN(n1205) );
  INVD1 U2797 ( .I(xi7_i[51]), .ZN(n1366) );
  INVD1 U2798 ( .I(xi7_r[51]), .ZN(n1236) );
  INVD1 U2799 ( .I(xi5_i[51]), .ZN(n1334) );
  INVD1 U2800 ( .I(xi5_r[51]), .ZN(n1204) );
  IND2D1 U2801 ( .A1(xi3_i[47]), .B1(xi7_i[47]), .ZN(sub_344_carry[1]) );
  INVD1 U2802 ( .I(xi7_i[48]), .ZN(n1369) );
  INVD1 U2803 ( .I(xi7_i[52]), .ZN(n1365) );
  IND2D1 U2804 ( .A1(xi3_r[47]), .B1(xi7_r[47]), .ZN(sub_335_carry[1]) );
  INVD1 U2805 ( .I(xi7_r[48]), .ZN(n1239) );
  INVD1 U2806 ( .I(xi7_r[52]), .ZN(n1235) );
  IND2D1 U2807 ( .A1(xi1_i[47]), .B1(xi5_i[47]), .ZN(sub_342_carry[1]) );
  INVD1 U2808 ( .I(xi5_i[48]), .ZN(n1337) );
  INVD1 U2809 ( .I(xi5_i[52]), .ZN(n1333) );
  IND2D1 U2810 ( .A1(xi1_r[47]), .B1(xi5_r[47]), .ZN(sub_333_carry[1]) );
  INVD1 U2811 ( .I(xi5_r[48]), .ZN(n1207) );
  INVD1 U2812 ( .I(xi5_r[52]), .ZN(n1203) );
  INVD1 U2813 ( .I(xi7_i[53]), .ZN(n1364) );
  INVD1 U2814 ( .I(xi7_r[53]), .ZN(n1234) );
  INVD1 U2815 ( .I(xi5_i[53]), .ZN(n1332) );
  INVD1 U2816 ( .I(xi5_r[53]), .ZN(n1202) );
  INVD1 U2817 ( .I(xi7_r[54]), .ZN(n1233) );
  INVD1 U2818 ( .I(xi5_r[54]), .ZN(n1201) );
  INVD1 U2819 ( .I(xi7_i[54]), .ZN(n1363) );
  INVD1 U2820 ( .I(xi7_r[55]), .ZN(n1232) );
  INVD1 U2821 ( .I(xi5_i[54]), .ZN(n1331) );
  INVD1 U2822 ( .I(xi5_r[55]), .ZN(n1200) );
  INVD1 U2823 ( .I(xi7_i[55]), .ZN(n1362) );
  INVD1 U2824 ( .I(xi7_r[56]), .ZN(n1231) );
  INVD1 U2825 ( .I(xi5_i[55]), .ZN(n1330) );
  INVD1 U2826 ( .I(xi5_r[56]), .ZN(n1199) );
  INVD1 U2827 ( .I(xi7_i[56]), .ZN(n1361) );
  INVD1 U2828 ( .I(xi7_r[57]), .ZN(n1230) );
  INVD1 U2829 ( .I(xi5_i[56]), .ZN(n1329) );
  INVD1 U2830 ( .I(xi5_r[57]), .ZN(n1198) );
  INVD1 U2831 ( .I(xi7_i[57]), .ZN(n1360) );
  INVD1 U2832 ( .I(xi7_r[58]), .ZN(n1229) );
  INVD1 U2833 ( .I(xi5_i[57]), .ZN(n1328) );
  INVD1 U2834 ( .I(xi5_r[58]), .ZN(n1197) );
  INVD1 U2835 ( .I(xi7_i[58]), .ZN(n1359) );
  INVD1 U2836 ( .I(xi7_r[59]), .ZN(n1228) );
  INVD1 U2837 ( .I(xi5_i[58]), .ZN(n1327) );
  INVD1 U2838 ( .I(xi5_r[59]), .ZN(n1196) );
  INVD1 U2839 ( .I(xi7_i[59]), .ZN(n1358) );
  INVD1 U2840 ( .I(xi7_r[60]), .ZN(n1227) );
  INVD1 U2841 ( .I(xi5_i[59]), .ZN(n1326) );
  INVD1 U2842 ( .I(xi5_r[60]), .ZN(n1195) );
  INVD1 U2843 ( .I(xi7_i[60]), .ZN(n1357) );
  INVD1 U2844 ( .I(xi7_r[61]), .ZN(n1226) );
  INVD1 U2845 ( .I(xi5_i[60]), .ZN(n1325) );
  INVD1 U2846 ( .I(xi5_r[61]), .ZN(n1194) );
  INVD1 U2847 ( .I(xi7_i[61]), .ZN(n1356) );
  INVD1 U2848 ( .I(xi7_r[62]), .ZN(n1225) );
  INVD1 U2849 ( .I(xi5_i[61]), .ZN(n1324) );
  INVD1 U2850 ( .I(xi5_r[62]), .ZN(n1193) );
  INVD1 U2851 ( .I(xi7_i[62]), .ZN(n1355) );
  INVD1 U2852 ( .I(xi5_i[62]), .ZN(n1323) );
  HA1D0 U2853 ( .A(dp_cluster_1_mult_512_C418_n246), .B(
        dp_cluster_1_mult_512_C418_n310), .CO(dp_cluster_1_mult_512_C418_n220), 
        .S(dp_cluster_1_mult_512_C418_n221) );
  OAI22D1 U2854 ( .A1(n2226), .A2(n976), .B1(n2304), .B2(n2225), .ZN(
        dp_cluster_1_mult_512_C418_n310) );
  OAI32D1 U2855 ( .A1(n1030), .A2(W3_8_i[48]), .A3(n2304), .B1(n1030), .B2(
        n976), .ZN(dp_cluster_1_mult_512_C418_n246) );
  HA1D0 U2856 ( .A(dp_cluster_1_mult_513_C418_n246), .B(
        dp_cluster_1_mult_513_C418_n310), .CO(dp_cluster_1_mult_513_C418_n220), 
        .S(dp_cluster_1_mult_513_C418_n221) );
  OAI22D1 U2857 ( .A1(n2074), .A2(n970), .B1(n2152), .B2(n2073), .ZN(
        dp_cluster_1_mult_513_C418_n310) );
  OAI32D1 U2858 ( .A1(n1074), .A2(W3_8_r[48]), .A3(n2152), .B1(n1074), .B2(
        n970), .ZN(dp_cluster_1_mult_513_C418_n246) );
  HA1D0 U2859 ( .A(dp_cluster_0_mult_485_C412_n246), .B(
        dp_cluster_0_mult_485_C412_n310), .CO(dp_cluster_0_mult_485_C412_n220), 
        .S(dp_cluster_0_mult_485_C412_n221) );
  OAI22D1 U2860 ( .A1(n1900), .A2(n964), .B1(n1978), .B2(n1899), .ZN(
        dp_cluster_0_mult_485_C412_n310) );
  OAI32D1 U2861 ( .A1(n1030), .A2(W3_8_r[48]), .A3(n1978), .B1(n1030), .B2(
        n964), .ZN(dp_cluster_0_mult_485_C412_n246) );
  HA1D0 U2862 ( .A(dp_cluster_3_mult_512_C415_n246), .B(
        dp_cluster_3_mult_512_C415_n310), .CO(dp_cluster_3_mult_512_C415_n220), 
        .S(dp_cluster_3_mult_512_C415_n221) );
  OAI22D1 U2863 ( .A1(n2877), .A2(n1000), .B1(n2955), .B2(n2876), .ZN(
        dp_cluster_3_mult_512_C415_n310) );
  OAI32D1 U2864 ( .A1(n1008), .A2(W1_8_i[48]), .A3(n2955), .B1(n1008), .B2(
        n1000), .ZN(dp_cluster_3_mult_512_C415_n246) );
  HA1D0 U2865 ( .A(dp_cluster_3_mult_513_C415_n246), .B(
        dp_cluster_3_mult_513_C415_n310), .CO(dp_cluster_3_mult_513_C415_n220), 
        .S(dp_cluster_3_mult_513_C415_n221) );
  OAI22D1 U2866 ( .A1(n2725), .A2(n994), .B1(n2803), .B2(n2724), .ZN(
        dp_cluster_3_mult_513_C415_n310) );
  OAI32D1 U2867 ( .A1(n1052), .A2(W1_8_r[48]), .A3(n2803), .B1(n1052), .B2(
        n994), .ZN(dp_cluster_3_mult_513_C415_n246) );
  HA1D0 U2868 ( .A(dp_cluster_2_mult_485_C409_n246), .B(
        dp_cluster_2_mult_485_C409_n310), .CO(dp_cluster_2_mult_485_C409_n220), 
        .S(dp_cluster_2_mult_485_C409_n221) );
  OAI22D1 U2869 ( .A1(n2551), .A2(n988), .B1(n2629), .B2(n2550), .ZN(
        dp_cluster_2_mult_485_C409_n310) );
  OAI32D1 U2870 ( .A1(n1008), .A2(W1_8_r[48]), .A3(n2629), .B1(n1008), .B2(
        n988), .ZN(dp_cluster_2_mult_485_C409_n246) );
  HA1D0 U2871 ( .A(dp_cluster_0_mult_486_C412_n246), .B(
        dp_cluster_0_mult_486_C412_n310), .CO(dp_cluster_0_mult_486_C412_n220), 
        .S(dp_cluster_0_mult_486_C412_n221) );
  OAI22D1 U2872 ( .A1(n1748), .A2(n958), .B1(n1826), .B2(n1747), .ZN(
        dp_cluster_0_mult_486_C412_n310) );
  OAI32D1 U2873 ( .A1(n1074), .A2(W3_8_i[48]), .A3(n1826), .B1(n1074), .B2(
        n958), .ZN(dp_cluster_0_mult_486_C412_n246) );
  HA1D0 U2874 ( .A(dp_cluster_2_mult_486_C409_n246), .B(
        dp_cluster_2_mult_486_C409_n310), .CO(dp_cluster_2_mult_486_C409_n220), 
        .S(dp_cluster_2_mult_486_C409_n221) );
  OAI22D1 U2875 ( .A1(n2399), .A2(n982), .B1(n2477), .B2(n2398), .ZN(
        dp_cluster_2_mult_486_C409_n310) );
  OAI32D1 U2876 ( .A1(n1052), .A2(W1_8_i[48]), .A3(n2477), .B1(n1052), .B2(
        n982), .ZN(dp_cluster_2_mult_486_C409_n246) );
  HA1D0 U2877 ( .A(dp_cluster_0_mult_485_C412_n248), .B(
        dp_cluster_0_mult_485_C412_n343), .CO(dp_cluster_0_mult_485_C412_n237), 
        .S(dp_cluster_0_mult_485_C412_n238) );
  OAI22D1 U2878 ( .A1(n1935), .A2(n960), .B1(n1936), .B2(n1933), .ZN(
        dp_cluster_0_mult_485_C412_n343) );
  OAI32D1 U2879 ( .A1(n1036), .A2(W3_8_r[48]), .A3(n1936), .B1(n1036), .B2(
        n960), .ZN(dp_cluster_0_mult_485_C412_n248) );
  HA1D0 U2880 ( .A(dp_cluster_2_mult_485_C409_n248), .B(
        dp_cluster_2_mult_485_C409_n343), .CO(dp_cluster_2_mult_485_C409_n237), 
        .S(dp_cluster_2_mult_485_C409_n238) );
  OAI22D1 U2881 ( .A1(n2586), .A2(n984), .B1(n2587), .B2(n2584), .ZN(
        dp_cluster_2_mult_485_C409_n343) );
  OAI32D1 U2882 ( .A1(n1014), .A2(W1_8_r[48]), .A3(n2587), .B1(n1014), .B2(
        n984), .ZN(dp_cluster_2_mult_485_C409_n248) );
  HA1D0 U2883 ( .A(dp_cluster_1_mult_513_C418_n248), .B(
        dp_cluster_1_mult_513_C418_n343), .CO(dp_cluster_1_mult_513_C418_n237), 
        .S(dp_cluster_1_mult_513_C418_n238) );
  OAI22D1 U2884 ( .A1(n2109), .A2(n966), .B1(n2110), .B2(n2107), .ZN(
        dp_cluster_1_mult_513_C418_n343) );
  OAI32D1 U2885 ( .A1(n1080), .A2(W3_8_r[48]), .A3(n2110), .B1(n1080), .B2(
        n966), .ZN(dp_cluster_1_mult_513_C418_n248) );
  HA1D0 U2886 ( .A(dp_cluster_3_mult_513_C415_n248), .B(
        dp_cluster_3_mult_513_C415_n343), .CO(dp_cluster_3_mult_513_C415_n237), 
        .S(dp_cluster_3_mult_513_C415_n238) );
  OAI22D1 U2887 ( .A1(n2760), .A2(n990), .B1(n2761), .B2(n2758), .ZN(
        dp_cluster_3_mult_513_C415_n343) );
  OAI32D1 U2888 ( .A1(n1058), .A2(W1_8_r[48]), .A3(n2761), .B1(n1058), .B2(
        n990), .ZN(dp_cluster_3_mult_513_C415_n248) );
  HA1D0 U2889 ( .A(dp_cluster_1_mult_512_C418_n248), .B(
        dp_cluster_1_mult_512_C418_n343), .CO(dp_cluster_1_mult_512_C418_n237), 
        .S(dp_cluster_1_mult_512_C418_n238) );
  OAI22D1 U2890 ( .A1(n2261), .A2(n972), .B1(n2262), .B2(n2259), .ZN(
        dp_cluster_1_mult_512_C418_n343) );
  OAI32D1 U2891 ( .A1(n1036), .A2(W3_8_i[48]), .A3(n2262), .B1(n1036), .B2(
        n972), .ZN(dp_cluster_1_mult_512_C418_n248) );
  HA1D0 U2892 ( .A(dp_cluster_3_mult_512_C415_n248), .B(
        dp_cluster_3_mult_512_C415_n343), .CO(dp_cluster_3_mult_512_C415_n237), 
        .S(dp_cluster_3_mult_512_C415_n238) );
  OAI22D1 U2893 ( .A1(n2912), .A2(n996), .B1(n2913), .B2(n2910), .ZN(
        dp_cluster_3_mult_512_C415_n343) );
  OAI32D1 U2894 ( .A1(n1014), .A2(W1_8_i[48]), .A3(n2913), .B1(n1014), .B2(
        n996), .ZN(dp_cluster_3_mult_512_C415_n248) );
  HA1D0 U2895 ( .A(dp_cluster_0_mult_486_C412_n248), .B(
        dp_cluster_0_mult_486_C412_n343), .CO(dp_cluster_0_mult_486_C412_n237), 
        .S(dp_cluster_0_mult_486_C412_n238) );
  OAI22D1 U2896 ( .A1(n1783), .A2(n954), .B1(n1784), .B2(n1781), .ZN(
        dp_cluster_0_mult_486_C412_n343) );
  OAI32D1 U2897 ( .A1(n1080), .A2(W3_8_i[48]), .A3(n1784), .B1(n1080), .B2(
        n954), .ZN(dp_cluster_0_mult_486_C412_n248) );
  HA1D0 U2898 ( .A(dp_cluster_2_mult_486_C409_n248), .B(
        dp_cluster_2_mult_486_C409_n343), .CO(dp_cluster_2_mult_486_C409_n237), 
        .S(dp_cluster_2_mult_486_C409_n238) );
  OAI22D1 U2899 ( .A1(n2434), .A2(n978), .B1(n2435), .B2(n2432), .ZN(
        dp_cluster_2_mult_486_C409_n343) );
  OAI32D1 U2900 ( .A1(n1058), .A2(W1_8_i[48]), .A3(n2435), .B1(n1058), .B2(
        n978), .ZN(dp_cluster_2_mult_486_C409_n248) );
  FA1D0 U2901 ( .A(dp_cluster_0_mult_485_C412_n242), .B(
        dp_cluster_0_mult_485_C412_n249), .CI(dp_cluster_0_mult_485_C412_n76), 
        .CO(dp_cluster_0_mult_485_C412_n75), .S(dp_cluster_0_N60) );
  OAI32D1 U2902 ( .A1(n1039), .A2(W3_8_r[48]), .A3(n1954), .B1(n1039), .B2(
        n961), .ZN(dp_cluster_0_mult_485_C412_n249) );
  FA1D0 U2903 ( .A(dp_cluster_2_mult_485_C409_n242), .B(
        dp_cluster_2_mult_485_C409_n249), .CI(dp_cluster_2_mult_485_C409_n76), 
        .CO(dp_cluster_2_mult_485_C409_n75), .S(dp_cluster_2_N4) );
  OAI32D1 U2904 ( .A1(n1017), .A2(W1_8_r[48]), .A3(n2605), .B1(n1017), .B2(
        n985), .ZN(dp_cluster_2_mult_485_C409_n249) );
  HA1D0 U2905 ( .A(dp_cluster_1_mult_512_C418_n244), .B(
        dp_cluster_1_mult_512_C418_n279), .CO(dp_cluster_1_mult_512_C418_n191), 
        .S(dp_cluster_1_mult_512_C418_n192) );
  OAI22D1 U2906 ( .A1(n2198), .A2(n975), .B1(n2310), .B2(n2197), .ZN(
        dp_cluster_1_mult_512_C418_n279) );
  OAI32D1 U2907 ( .A1(n1025), .A2(W3_8_i[48]), .A3(n2310), .B1(n1025), .B2(
        n975), .ZN(dp_cluster_1_mult_512_C418_n244) );
  HA1D0 U2908 ( .A(dp_cluster_1_mult_513_C418_n244), .B(
        dp_cluster_1_mult_513_C418_n279), .CO(dp_cluster_1_mult_513_C418_n191), 
        .S(dp_cluster_1_mult_513_C418_n192) );
  OAI22D1 U2909 ( .A1(n2046), .A2(n969), .B1(n2158), .B2(n2045), .ZN(
        dp_cluster_1_mult_513_C418_n279) );
  OAI32D1 U2910 ( .A1(n1069), .A2(W3_8_r[48]), .A3(n2158), .B1(n1069), .B2(
        n969), .ZN(dp_cluster_1_mult_513_C418_n244) );
  HA1D0 U2911 ( .A(dp_cluster_0_mult_486_C412_n244), .B(
        dp_cluster_0_mult_486_C412_n279), .CO(dp_cluster_0_mult_486_C412_n191), 
        .S(dp_cluster_0_mult_486_C412_n192) );
  OAI22D1 U2912 ( .A1(n1720), .A2(n957), .B1(n1832), .B2(n1719), .ZN(
        dp_cluster_0_mult_486_C412_n279) );
  OAI32D1 U2913 ( .A1(n1069), .A2(W3_8_i[48]), .A3(n1832), .B1(n1069), .B2(
        n957), .ZN(dp_cluster_0_mult_486_C412_n244) );
  HA1D0 U2914 ( .A(dp_cluster_0_mult_485_C412_n244), .B(
        dp_cluster_0_mult_485_C412_n279), .CO(dp_cluster_0_mult_485_C412_n191), 
        .S(dp_cluster_0_mult_485_C412_n192) );
  OAI22D1 U2915 ( .A1(n1872), .A2(n963), .B1(n1984), .B2(n1871), .ZN(
        dp_cluster_0_mult_485_C412_n279) );
  OAI32D1 U2916 ( .A1(n1025), .A2(W3_8_r[48]), .A3(n1984), .B1(n1025), .B2(
        n963), .ZN(dp_cluster_0_mult_485_C412_n244) );
  HA1D0 U2917 ( .A(dp_cluster_3_mult_512_C415_n244), .B(
        dp_cluster_3_mult_512_C415_n279), .CO(dp_cluster_3_mult_512_C415_n191), 
        .S(dp_cluster_3_mult_512_C415_n192) );
  OAI22D1 U2918 ( .A1(n2849), .A2(n999), .B1(n2961), .B2(n2848), .ZN(
        dp_cluster_3_mult_512_C415_n279) );
  OAI32D1 U2919 ( .A1(n1003), .A2(W1_8_i[48]), .A3(n2961), .B1(n1003), .B2(
        n999), .ZN(dp_cluster_3_mult_512_C415_n244) );
  HA1D0 U2920 ( .A(dp_cluster_3_mult_513_C415_n244), .B(
        dp_cluster_3_mult_513_C415_n279), .CO(dp_cluster_3_mult_513_C415_n191), 
        .S(dp_cluster_3_mult_513_C415_n192) );
  OAI22D1 U2921 ( .A1(n2697), .A2(n993), .B1(n2809), .B2(n2696), .ZN(
        dp_cluster_3_mult_513_C415_n279) );
  OAI32D1 U2922 ( .A1(n1047), .A2(W1_8_r[48]), .A3(n2809), .B1(n1047), .B2(
        n993), .ZN(dp_cluster_3_mult_513_C415_n244) );
  HA1D0 U2923 ( .A(dp_cluster_2_mult_486_C409_n244), .B(
        dp_cluster_2_mult_486_C409_n279), .CO(dp_cluster_2_mult_486_C409_n191), 
        .S(dp_cluster_2_mult_486_C409_n192) );
  OAI22D1 U2924 ( .A1(n2371), .A2(n981), .B1(n2483), .B2(n2370), .ZN(
        dp_cluster_2_mult_486_C409_n279) );
  OAI32D1 U2925 ( .A1(n1047), .A2(W1_8_i[48]), .A3(n2483), .B1(n1047), .B2(
        n981), .ZN(dp_cluster_2_mult_486_C409_n244) );
  HA1D0 U2926 ( .A(dp_cluster_2_mult_485_C409_n244), .B(
        dp_cluster_2_mult_485_C409_n279), .CO(dp_cluster_2_mult_485_C409_n191), 
        .S(dp_cluster_2_mult_485_C409_n192) );
  OAI22D1 U2927 ( .A1(n2523), .A2(n987), .B1(n2635), .B2(n2522), .ZN(
        dp_cluster_2_mult_485_C409_n279) );
  OAI32D1 U2928 ( .A1(n1003), .A2(W1_8_r[48]), .A3(n2635), .B1(n1003), .B2(
        n987), .ZN(dp_cluster_2_mult_485_C409_n244) );
  HA1D0 U2929 ( .A(dp_cluster_1_mult_513_C418_n247), .B(
        dp_cluster_1_mult_513_C418_n327), .CO(dp_cluster_1_mult_513_C418_n230), 
        .S(dp_cluster_1_mult_513_C418_n231) );
  OAI22D1 U2930 ( .A1(n2091), .A2(n968), .B1(n2092), .B2(n2089), .ZN(
        dp_cluster_1_mult_513_C418_n327) );
  OAI32D1 U2931 ( .A1(n1077), .A2(W3_8_r[48]), .A3(n2092), .B1(n1077), .B2(
        n968), .ZN(dp_cluster_1_mult_513_C418_n247) );
  HA1D0 U2932 ( .A(dp_cluster_3_mult_513_C415_n247), .B(
        dp_cluster_3_mult_513_C415_n327), .CO(dp_cluster_3_mult_513_C415_n230), 
        .S(dp_cluster_3_mult_513_C415_n231) );
  OAI22D1 U2933 ( .A1(n2742), .A2(n992), .B1(n2743), .B2(n2740), .ZN(
        dp_cluster_3_mult_513_C415_n327) );
  OAI32D1 U2934 ( .A1(n1055), .A2(W1_8_r[48]), .A3(n2743), .B1(n1055), .B2(
        n992), .ZN(dp_cluster_3_mult_513_C415_n247) );
  HA1D0 U2935 ( .A(dp_cluster_1_mult_512_C418_n247), .B(
        dp_cluster_1_mult_512_C418_n327), .CO(dp_cluster_1_mult_512_C418_n230), 
        .S(dp_cluster_1_mult_512_C418_n231) );
  OAI22D1 U2936 ( .A1(n2243), .A2(n974), .B1(n2244), .B2(n2241), .ZN(
        dp_cluster_1_mult_512_C418_n327) );
  OAI32D1 U2937 ( .A1(n1033), .A2(W3_8_i[48]), .A3(n2244), .B1(n1033), .B2(
        n974), .ZN(dp_cluster_1_mult_512_C418_n247) );
  HA1D0 U2938 ( .A(dp_cluster_3_mult_512_C415_n247), .B(
        dp_cluster_3_mult_512_C415_n327), .CO(dp_cluster_3_mult_512_C415_n230), 
        .S(dp_cluster_3_mult_512_C415_n231) );
  OAI22D1 U2939 ( .A1(n2894), .A2(n998), .B1(n2895), .B2(n2892), .ZN(
        dp_cluster_3_mult_512_C415_n327) );
  OAI32D1 U2940 ( .A1(n1011), .A2(W1_8_i[48]), .A3(n2895), .B1(n1011), .B2(
        n998), .ZN(dp_cluster_3_mult_512_C415_n247) );
  HA1D0 U2941 ( .A(dp_cluster_0_mult_486_C412_n243), .B(
        dp_cluster_0_mult_486_C412_n263), .CO(dp_cluster_0_mult_486_C412_n172), 
        .S(dp_cluster_0_mult_486_C412_n173) );
  OAI22D1 U2942 ( .A1(n1706), .A2(n1828), .B1(n1829), .B2(n1705), .ZN(
        dp_cluster_0_mult_486_C412_n263) );
  OAI32D1 U2943 ( .A1(n1067), .A2(W3_8_i[48]), .A3(n1829), .B1(n1067), .B2(
        n1828), .ZN(dp_cluster_0_mult_486_C412_n243) );
  HA1D0 U2944 ( .A(dp_cluster_0_mult_485_C412_n243), .B(
        dp_cluster_0_mult_485_C412_n263), .CO(dp_cluster_0_mult_485_C412_n172), 
        .S(dp_cluster_0_mult_485_C412_n173) );
  OAI22D1 U2945 ( .A1(n1858), .A2(n1980), .B1(n1981), .B2(n1857), .ZN(
        dp_cluster_0_mult_485_C412_n263) );
  OAI32D1 U2946 ( .A1(n1023), .A2(W3_8_r[48]), .A3(n1981), .B1(n1023), .B2(
        n1980), .ZN(dp_cluster_0_mult_485_C412_n243) );
  HA1D0 U2947 ( .A(dp_cluster_2_mult_486_C409_n243), .B(
        dp_cluster_2_mult_486_C409_n263), .CO(dp_cluster_2_mult_486_C409_n172), 
        .S(dp_cluster_2_mult_486_C409_n173) );
  OAI22D1 U2948 ( .A1(n2357), .A2(n2479), .B1(n2480), .B2(n2356), .ZN(
        dp_cluster_2_mult_486_C409_n263) );
  OAI32D1 U2949 ( .A1(n1045), .A2(W1_8_i[48]), .A3(n2480), .B1(n1045), .B2(
        n2479), .ZN(dp_cluster_2_mult_486_C409_n243) );
  HA1D0 U2950 ( .A(dp_cluster_2_mult_485_C409_n243), .B(
        dp_cluster_2_mult_485_C409_n263), .CO(dp_cluster_2_mult_485_C409_n172), 
        .S(dp_cluster_2_mult_485_C409_n173) );
  OAI22D1 U2951 ( .A1(n2509), .A2(n2631), .B1(n2632), .B2(n2508), .ZN(
        dp_cluster_2_mult_485_C409_n263) );
  OAI32D1 U2952 ( .A1(n1001), .A2(W1_8_r[48]), .A3(n2632), .B1(n1001), .B2(
        n2631), .ZN(dp_cluster_2_mult_485_C409_n243) );
  HA1D0 U2953 ( .A(dp_cluster_1_mult_512_C418_n245), .B(
        dp_cluster_1_mult_512_C418_n294), .CO(dp_cluster_1_mult_512_C418_n207), 
        .S(dp_cluster_1_mult_512_C418_n208) );
  OAI22D1 U2954 ( .A1(n2212), .A2(n971), .B1(n2300), .B2(n2211), .ZN(
        dp_cluster_1_mult_512_C418_n294) );
  OAI32D1 U2955 ( .A1(n1028), .A2(W3_8_i[48]), .A3(n2300), .B1(n1028), .B2(
        n971), .ZN(dp_cluster_1_mult_512_C418_n245) );
  HA1D0 U2956 ( .A(dp_cluster_1_mult_513_C418_n245), .B(
        dp_cluster_1_mult_513_C418_n294), .CO(dp_cluster_1_mult_513_C418_n207), 
        .S(dp_cluster_1_mult_513_C418_n208) );
  OAI22D1 U2957 ( .A1(n2060), .A2(n965), .B1(n2148), .B2(n2059), .ZN(
        dp_cluster_1_mult_513_C418_n294) );
  OAI32D1 U2958 ( .A1(n1072), .A2(W3_8_r[48]), .A3(n2148), .B1(n1072), .B2(
        n965), .ZN(dp_cluster_1_mult_513_C418_n245) );
  HA1D0 U2959 ( .A(dp_cluster_0_mult_486_C412_n245), .B(
        dp_cluster_0_mult_486_C412_n294), .CO(dp_cluster_0_mult_486_C412_n207), 
        .S(dp_cluster_0_mult_486_C412_n208) );
  OAI22D1 U2960 ( .A1(n1734), .A2(n953), .B1(n1822), .B2(n1733), .ZN(
        dp_cluster_0_mult_486_C412_n294) );
  OAI32D1 U2961 ( .A1(n1072), .A2(W3_8_i[48]), .A3(n1822), .B1(n1072), .B2(
        n953), .ZN(dp_cluster_0_mult_486_C412_n245) );
  HA1D0 U2962 ( .A(dp_cluster_0_mult_485_C412_n245), .B(
        dp_cluster_0_mult_485_C412_n294), .CO(dp_cluster_0_mult_485_C412_n207), 
        .S(dp_cluster_0_mult_485_C412_n208) );
  OAI22D1 U2963 ( .A1(n1886), .A2(n959), .B1(n1974), .B2(n1885), .ZN(
        dp_cluster_0_mult_485_C412_n294) );
  OAI32D1 U2964 ( .A1(n1028), .A2(W3_8_r[48]), .A3(n1974), .B1(n1028), .B2(
        n959), .ZN(dp_cluster_0_mult_485_C412_n245) );
  HA1D0 U2965 ( .A(dp_cluster_3_mult_512_C415_n245), .B(
        dp_cluster_3_mult_512_C415_n294), .CO(dp_cluster_3_mult_512_C415_n207), 
        .S(dp_cluster_3_mult_512_C415_n208) );
  OAI22D1 U2966 ( .A1(n2863), .A2(n995), .B1(n2951), .B2(n2862), .ZN(
        dp_cluster_3_mult_512_C415_n294) );
  OAI32D1 U2967 ( .A1(n1006), .A2(W1_8_i[48]), .A3(n2951), .B1(n1006), .B2(
        n995), .ZN(dp_cluster_3_mult_512_C415_n245) );
  HA1D0 U2968 ( .A(dp_cluster_3_mult_513_C415_n245), .B(
        dp_cluster_3_mult_513_C415_n294), .CO(dp_cluster_3_mult_513_C415_n207), 
        .S(dp_cluster_3_mult_513_C415_n208) );
  OAI22D1 U2969 ( .A1(n2711), .A2(n989), .B1(n2799), .B2(n2710), .ZN(
        dp_cluster_3_mult_513_C415_n294) );
  OAI32D1 U2970 ( .A1(n1050), .A2(W1_8_r[48]), .A3(n2799), .B1(n1050), .B2(
        n989), .ZN(dp_cluster_3_mult_513_C415_n245) );
  HA1D0 U2971 ( .A(dp_cluster_2_mult_486_C409_n245), .B(
        dp_cluster_2_mult_486_C409_n294), .CO(dp_cluster_2_mult_486_C409_n207), 
        .S(dp_cluster_2_mult_486_C409_n208) );
  OAI22D1 U2972 ( .A1(n2385), .A2(n977), .B1(n2473), .B2(n2384), .ZN(
        dp_cluster_2_mult_486_C409_n294) );
  OAI32D1 U2973 ( .A1(n1050), .A2(W1_8_i[48]), .A3(n2473), .B1(n1050), .B2(
        n977), .ZN(dp_cluster_2_mult_486_C409_n245) );
  HA1D0 U2974 ( .A(dp_cluster_2_mult_485_C409_n245), .B(
        dp_cluster_2_mult_485_C409_n294), .CO(dp_cluster_2_mult_485_C409_n207), 
        .S(dp_cluster_2_mult_485_C409_n208) );
  OAI22D1 U2975 ( .A1(n2537), .A2(n983), .B1(n2625), .B2(n2536), .ZN(
        dp_cluster_2_mult_485_C409_n294) );
  OAI32D1 U2976 ( .A1(n1006), .A2(W1_8_r[48]), .A3(n2625), .B1(n1006), .B2(
        n983), .ZN(dp_cluster_2_mult_485_C409_n245) );
  HA1D0 U2977 ( .A(dp_cluster_0_mult_485_C412_n376), .B(
        dp_cluster_0_mult_485_C412_n250), .CO(dp_cluster_0_mult_485_C412_n77), 
        .S(dp_cluster_0_N58) );
  IOA21D1 U2978 ( .A1(n1094), .A2(n1109), .B(n1970), .ZN(
        dp_cluster_0_mult_485_C412_n250) );
  OAI22D1 U2979 ( .A1(W3_8_r[48]), .A2(n1970), .B1(n1969), .B2(n1043), .ZN(
        dp_cluster_0_mult_485_C412_n376) );
  HA1D0 U2980 ( .A(dp_cluster_2_mult_485_C409_n376), .B(
        dp_cluster_2_mult_485_C409_n250), .CO(dp_cluster_2_mult_485_C409_n77), 
        .S(dp_cluster_2_N2) );
  IOA21D1 U2981 ( .A1(n1091), .A2(n1112), .B(n2621), .ZN(
        dp_cluster_2_mult_485_C409_n250) );
  OAI22D1 U2982 ( .A1(W1_8_r[48]), .A2(n2621), .B1(n2620), .B2(n1021), .ZN(
        dp_cluster_2_mult_485_C409_n376) );
  INVD1 U2983 ( .I(W3_8_i[48]), .ZN(n1429) );
  INVD1 U2984 ( .I(W1_8_i[48]), .ZN(n1414) );
  OAI22D1 U2985 ( .A1(n2312), .A2(n975), .B1(n2310), .B2(n2309), .ZN(n2313) );
  OAI22D1 U2986 ( .A1(n2963), .A2(n999), .B1(n2961), .B2(n2960), .ZN(n2964) );
  INVD1 U2987 ( .I(xo2_i_w_d1r[14]), .ZN(n1527) );
  INVD1 U2988 ( .I(xo2_r_w_d1r[14]), .ZN(n1511) );
  INVD1 U2989 ( .I(xo6_r_w_d1r[14]), .ZN(n1639) );
  INVD1 U2990 ( .I(xo6_i_w_d1r[14]), .ZN(n1655) );
  INVD1 U2991 ( .I(xo2_i_w_d1r[15]), .ZN(n1526) );
  INVD1 U2992 ( .I(xo2_r_w_d1r[15]), .ZN(n1510) );
  INVD1 U2993 ( .I(xo6_r_w_d1r[15]), .ZN(n1638) );
  INVD1 U2994 ( .I(xo6_i_w_d1r[15]), .ZN(n1654) );
  INVD1 U2995 ( .I(xo3_i_w_d1r[3]), .ZN(n1554) );
  INVD1 U2996 ( .I(xo7_i_w_d1r[3]), .ZN(n1682) );
  INVD1 U2997 ( .I(xo1_r_w_d1r[14]), .ZN(n1435) );
  INVD1 U2998 ( .I(xo3_i_w_d1r[14]), .ZN(n1543) );
  INVD1 U2999 ( .I(xo1_r_w_d1r[15]), .ZN(n1432) );
  INVD1 U3000 ( .I(xo3_i_w_d1r[15]), .ZN(n1542) );
  INVD1 U3001 ( .I(xo7_i_w_d1r[14]), .ZN(n1671) );
  INVD1 U3002 ( .I(xo5_r_w_d1r[14]), .ZN(n1563) );
  INVD1 U3003 ( .I(xo5_r_w_d1r[15]), .ZN(n1560) );
  INVD1 U3004 ( .I(xo7_i_w_d1r[15]), .ZN(n1670) );
  INVD1 U3005 ( .I(xi6_r[49]), .ZN(n1222) );
  INVD1 U3006 ( .I(xi6_r[50]), .ZN(n1221) );
  INVD1 U3007 ( .I(xi6_r[51]), .ZN(n1220) );
  INVD1 U3008 ( .I(xi6_r[52]), .ZN(n1219) );
  INVD1 U3009 ( .I(xi6_r[53]), .ZN(n1218) );
  INVD1 U3010 ( .I(xi6_r[54]), .ZN(n1217) );
  INVD1 U3011 ( .I(xi6_r[55]), .ZN(n1216) );
  INVD1 U3012 ( .I(xi6_r[56]), .ZN(n1215) );
  INVD1 U3013 ( .I(xo1_r_w_d1r[2]), .ZN(n1471) );
  INVD1 U3014 ( .I(xo3_i_w_d1r[2]), .ZN(n1555) );
  ND2D1 U3015 ( .A1(xo2_i_w_d1r[0]), .A2(n949), .ZN(sub_360_carry[1]) );
  INVD1 U3016 ( .I(xo2_i_w_d1r[1]), .ZN(n1540) );
  INVD1 U3017 ( .I(xo0_i_w_d1r[0]), .ZN(n949) );
  ND2D1 U3018 ( .A1(xo2_r_w_d1r[0]), .A2(n951), .ZN(sub_351_carry[1]) );
  INVD1 U3019 ( .I(xo2_r_w_d1r[1]), .ZN(n1524) );
  INVD1 U3020 ( .I(xo0_r_w_d1r[0]), .ZN(n951) );
  ND2D1 U3021 ( .A1(xo6_r_w_d1r[0]), .A2(n950), .ZN(sub_355_carry[1]) );
  INVD1 U3022 ( .I(xo6_r_w_d1r[1]), .ZN(n1652) );
  INVD1 U3023 ( .I(xo4_r_w_d1r[0]), .ZN(n950) );
  ND2D1 U3024 ( .A1(xo6_i_w_d1r[0]), .A2(n947), .ZN(sub_364_carry[1]) );
  INVD1 U3025 ( .I(xo6_i_w_d1r[1]), .ZN(n1668) );
  INVD1 U3026 ( .I(xo4_i_w_d1r[0]), .ZN(n947) );
  INVD1 U3027 ( .I(xo1_r_w_d1r[3]), .ZN(n1468) );
  INVD1 U3028 ( .I(xo2_i_w_d1r[2]), .ZN(n1539) );
  INVD1 U3029 ( .I(xo2_r_w_d1r[2]), .ZN(n1523) );
  INVD1 U3030 ( .I(xo6_r_w_d1r[2]), .ZN(n1651) );
  INVD1 U3031 ( .I(xo7_i_w_d1r[2]), .ZN(n1683) );
  INVD1 U3032 ( .I(xo6_i_w_d1r[2]), .ZN(n1667) );
  INVD1 U3033 ( .I(xo5_r_w_d1r[2]), .ZN(n1599) );
  INVD1 U3034 ( .I(xi6_r[57]), .ZN(n1214) );
  INVD1 U3035 ( .I(xo1_r_w_d1r[4]), .ZN(n1465) );
  INVD1 U3036 ( .I(xo3_i_w_d1r[4]), .ZN(n1553) );
  INVD1 U3037 ( .I(xo2_i_w_d1r[3]), .ZN(n1538) );
  INVD1 U3038 ( .I(xo2_r_w_d1r[3]), .ZN(n1522) );
  INVD1 U3039 ( .I(xo6_r_w_d1r[3]), .ZN(n1650) );
  INVD1 U3040 ( .I(xo6_i_w_d1r[3]), .ZN(n1666) );
  INVD1 U3041 ( .I(xo5_r_w_d1r[3]), .ZN(n1596) );
  INVD1 U3042 ( .I(xo1_r_w_d1r[5]), .ZN(n1462) );
  INVD1 U3043 ( .I(xo3_i_w_d1r[5]), .ZN(n1552) );
  INVD1 U3044 ( .I(xo2_i_w_d1r[4]), .ZN(n1537) );
  INVD1 U3045 ( .I(xo2_r_w_d1r[4]), .ZN(n1521) );
  INVD1 U3046 ( .I(xo6_r_w_d1r[4]), .ZN(n1649) );
  INVD1 U3047 ( .I(xo7_i_w_d1r[4]), .ZN(n1681) );
  INVD1 U3048 ( .I(xo6_i_w_d1r[4]), .ZN(n1665) );
  INVD1 U3049 ( .I(xo5_r_w_d1r[4]), .ZN(n1593) );
  INVD1 U3050 ( .I(xi6_r[58]), .ZN(n1213) );
  INVD1 U3051 ( .I(xo1_r_w_d1r[6]), .ZN(n1459) );
  INVD1 U3052 ( .I(xo3_i_w_d1r[6]), .ZN(n1551) );
  INVD1 U3053 ( .I(xo2_i_w_d1r[5]), .ZN(n1536) );
  INVD1 U3054 ( .I(xo2_r_w_d1r[5]), .ZN(n1520) );
  INVD1 U3055 ( .I(xo6_r_w_d1r[5]), .ZN(n1648) );
  INVD1 U3056 ( .I(xo7_i_w_d1r[5]), .ZN(n1680) );
  INVD1 U3057 ( .I(xo6_i_w_d1r[5]), .ZN(n1664) );
  INVD1 U3058 ( .I(xo5_r_w_d1r[5]), .ZN(n1590) );
  INVD1 U3059 ( .I(xo1_r_w_d1r[7]), .ZN(n1456) );
  INVD1 U3060 ( .I(xo3_i_w_d1r[7]), .ZN(n1550) );
  INVD1 U3061 ( .I(xo2_i_w_d1r[6]), .ZN(n1535) );
  INVD1 U3062 ( .I(xo2_r_w_d1r[6]), .ZN(n1519) );
  INVD1 U3063 ( .I(xo6_r_w_d1r[6]), .ZN(n1647) );
  INVD1 U3064 ( .I(xo7_i_w_d1r[6]), .ZN(n1679) );
  INVD1 U3065 ( .I(xo6_i_w_d1r[6]), .ZN(n1663) );
  INVD1 U3066 ( .I(xo5_r_w_d1r[6]), .ZN(n1587) );
  INVD1 U3067 ( .I(xi6_r[59]), .ZN(n1212) );
  INVD1 U3068 ( .I(xo1_r_w_d1r[8]), .ZN(n1453) );
  INVD1 U3069 ( .I(xo3_i_w_d1r[8]), .ZN(n1549) );
  INVD1 U3070 ( .I(xo2_i_w_d1r[7]), .ZN(n1534) );
  INVD1 U3071 ( .I(xo2_r_w_d1r[7]), .ZN(n1518) );
  INVD1 U3072 ( .I(xo6_r_w_d1r[7]), .ZN(n1646) );
  INVD1 U3073 ( .I(xo7_i_w_d1r[7]), .ZN(n1678) );
  INVD1 U3074 ( .I(xo6_i_w_d1r[7]), .ZN(n1662) );
  INVD1 U3075 ( .I(xo5_r_w_d1r[7]), .ZN(n1584) );
  INVD1 U3076 ( .I(xo1_r_w_d1r[9]), .ZN(n1450) );
  INVD1 U3077 ( .I(xo3_i_w_d1r[9]), .ZN(n1548) );
  INVD1 U3078 ( .I(xo2_i_w_d1r[8]), .ZN(n1533) );
  INVD1 U3079 ( .I(xo2_r_w_d1r[8]), .ZN(n1517) );
  INVD1 U3080 ( .I(xo6_r_w_d1r[8]), .ZN(n1645) );
  INVD1 U3081 ( .I(xo7_i_w_d1r[8]), .ZN(n1677) );
  INVD1 U3082 ( .I(xo6_i_w_d1r[8]), .ZN(n1661) );
  INVD1 U3083 ( .I(xo5_r_w_d1r[8]), .ZN(n1581) );
  INVD1 U3084 ( .I(xi6_r[60]), .ZN(n1211) );
  INVD1 U3085 ( .I(xo1_r_w_d1r[10]), .ZN(n1447) );
  INVD1 U3086 ( .I(xo3_i_w_d1r[10]), .ZN(n1547) );
  INVD1 U3087 ( .I(xo2_i_w_d1r[9]), .ZN(n1532) );
  INVD1 U3088 ( .I(xo2_r_w_d1r[9]), .ZN(n1516) );
  INVD1 U3089 ( .I(xo6_r_w_d1r[9]), .ZN(n1644) );
  INVD1 U3090 ( .I(xo7_i_w_d1r[9]), .ZN(n1676) );
  INVD1 U3091 ( .I(xo6_i_w_d1r[9]), .ZN(n1660) );
  INVD1 U3092 ( .I(xo5_r_w_d1r[9]), .ZN(n1578) );
  INVD1 U3093 ( .I(xo1_r_w_d1r[11]), .ZN(n1444) );
  INVD1 U3094 ( .I(xo3_i_w_d1r[11]), .ZN(n1546) );
  INVD1 U3095 ( .I(xo2_i_w_d1r[10]), .ZN(n1531) );
  INVD1 U3096 ( .I(xo2_r_w_d1r[10]), .ZN(n1515) );
  INVD1 U3097 ( .I(xo6_r_w_d1r[10]), .ZN(n1643) );
  INVD1 U3098 ( .I(xo7_i_w_d1r[10]), .ZN(n1675) );
  INVD1 U3099 ( .I(xo6_i_w_d1r[10]), .ZN(n1659) );
  INVD1 U3100 ( .I(xo5_r_w_d1r[10]), .ZN(n1575) );
  INVD1 U3101 ( .I(xi6_r[61]), .ZN(n1210) );
  INVD1 U3102 ( .I(xo1_r_w_d1r[12]), .ZN(n1441) );
  INVD1 U3103 ( .I(xo3_i_w_d1r[12]), .ZN(n1545) );
  INVD1 U3104 ( .I(xo2_i_w_d1r[11]), .ZN(n1530) );
  INVD1 U3105 ( .I(xo2_r_w_d1r[11]), .ZN(n1514) );
  INVD1 U3106 ( .I(xo6_r_w_d1r[11]), .ZN(n1642) );
  INVD1 U3107 ( .I(xo7_i_w_d1r[11]), .ZN(n1674) );
  INVD1 U3108 ( .I(xo6_i_w_d1r[11]), .ZN(n1658) );
  INVD1 U3109 ( .I(xo5_r_w_d1r[11]), .ZN(n1572) );
  INVD1 U3110 ( .I(xo1_r_w_d1r[13]), .ZN(n1438) );
  INVD1 U3111 ( .I(xo3_i_w_d1r[13]), .ZN(n1544) );
  INVD1 U3112 ( .I(xo2_i_w_d1r[12]), .ZN(n1529) );
  INVD1 U3113 ( .I(xo2_r_w_d1r[12]), .ZN(n1513) );
  INVD1 U3114 ( .I(xo6_r_w_d1r[12]), .ZN(n1641) );
  INVD1 U3115 ( .I(xo7_i_w_d1r[12]), .ZN(n1673) );
  INVD1 U3116 ( .I(xo6_i_w_d1r[12]), .ZN(n1657) );
  INVD1 U3117 ( .I(xo5_r_w_d1r[12]), .ZN(n1569) );
  INVD1 U3118 ( .I(xi6_r[62]), .ZN(n1209) );
  INVD1 U3119 ( .I(xo2_i_w_d1r[13]), .ZN(n1528) );
  INVD1 U3120 ( .I(xo2_r_w_d1r[13]), .ZN(n1512) );
  INVD1 U3121 ( .I(xo6_r_w_d1r[13]), .ZN(n1640) );
  INVD1 U3122 ( .I(xo7_i_w_d1r[13]), .ZN(n1672) );
  INVD1 U3123 ( .I(xo6_i_w_d1r[13]), .ZN(n1656) );
  INVD1 U3124 ( .I(xo5_r_w_d1r[13]), .ZN(n1566) );
  ND2D1 U3125 ( .A1(xo1_r_w_d1r[0]), .A2(n936), .ZN(
        dp_cluster_5_sub_1_root_sub_440_carry[1]) );
  INVD1 U3126 ( .I(xo1_r_w_d1r[1]), .ZN(n1474) );
  INVD1 U3127 ( .I(xo3_r_w_d1r[0]), .ZN(n936) );
  ND2D1 U3128 ( .A1(xo3_i_w_d1r[0]), .A2(n948), .ZN(sub_361_carry[1]) );
  INVD1 U3129 ( .I(xo3_i_w_d1r[1]), .ZN(n1556) );
  INVD1 U3130 ( .I(xo1_i_w_d1r[0]), .ZN(n948) );
  ND2D1 U3131 ( .A1(xo7_i_w_d1r[0]), .A2(n946), .ZN(sub_365_carry[1]) );
  INVD1 U3132 ( .I(xo7_i_w_d1r[1]), .ZN(n1684) );
  INVD1 U3133 ( .I(xo5_i_w_d1r[0]), .ZN(n946) );
  ND2D1 U3134 ( .A1(xo5_r_w_d1r[0]), .A2(n937), .ZN(
        dp_cluster_4_sub_1_root_sub_444_carry[1]) );
  INVD1 U3135 ( .I(xo5_r_w_d1r[1]), .ZN(n1602) );
  INVD1 U3136 ( .I(xo7_r_w_d1r[0]), .ZN(n937) );
  IND2D1 U3137 ( .A1(xi2_r[47]), .B1(xi6_r[47]), .ZN(sub_334_carry[1]) );
  INVD1 U3138 ( .I(xi6_r[48]), .ZN(n1223) );
  IND2D1 U3139 ( .A1(xi2_i[47]), .B1(xi6_i[47]), .ZN(sub_343_carry[1]) );
  INVD1 U3140 ( .I(xi6_i[48]), .ZN(n1353) );
  INVD1 U3141 ( .I(xi6_i[49]), .ZN(n1352) );
  INVD1 U3142 ( .I(xi6_i[50]), .ZN(n1351) );
  INVD1 U3143 ( .I(xi6_i[51]), .ZN(n1350) );
  INVD1 U3144 ( .I(xi6_i[52]), .ZN(n1349) );
  INVD1 U3145 ( .I(xi6_i[53]), .ZN(n1348) );
  INVD1 U3146 ( .I(xi6_i[54]), .ZN(n1347) );
  INVD1 U3147 ( .I(xi6_i[55]), .ZN(n1346) );
  INVD1 U3148 ( .I(xi6_i[56]), .ZN(n1345) );
  INVD1 U3149 ( .I(xi6_i[57]), .ZN(n1344) );
  INVD1 U3150 ( .I(xi6_i[58]), .ZN(n1343) );
  INVD1 U3151 ( .I(xi6_i[59]), .ZN(n1342) );
  INVD1 U3152 ( .I(xi6_i[60]), .ZN(n1341) );
  INVD1 U3153 ( .I(xi6_i[61]), .ZN(n1340) );
  INVD1 U3154 ( .I(xi6_i[62]), .ZN(n1339) );
  IND2D1 U3155 ( .A1(xi0_i[47]), .B1(xi4_i[47]), .ZN(sub_341_carry[1]) );
  INVD1 U3156 ( .I(xi4_i[48]), .ZN(n1321) );
  INVD1 U3157 ( .I(xi4_i[49]), .ZN(n1320) );
  INVD1 U3158 ( .I(xi4_i[50]), .ZN(n1319) );
  INVD1 U3159 ( .I(xi4_i[51]), .ZN(n1318) );
  INVD1 U3160 ( .I(xi4_i[52]), .ZN(n1317) );
  INVD1 U3161 ( .I(xi4_i[53]), .ZN(n1316) );
  INVD1 U3162 ( .I(xi4_i[54]), .ZN(n1315) );
  INVD1 U3163 ( .I(xi4_i[55]), .ZN(n1314) );
  INVD1 U3164 ( .I(xi4_i[56]), .ZN(n1313) );
  INVD1 U3165 ( .I(xi4_i[57]), .ZN(n1312) );
  INVD1 U3166 ( .I(xi4_i[58]), .ZN(n1311) );
  INVD1 U3167 ( .I(xi4_i[59]), .ZN(n1310) );
  INVD1 U3168 ( .I(xi4_i[60]), .ZN(n1309) );
  INVD1 U3169 ( .I(xi4_i[61]), .ZN(n1308) );
  INVD1 U3170 ( .I(xi4_i[62]), .ZN(n1307) );
  IND2D1 U3171 ( .A1(xi0_r[47]), .B1(xi4_r[47]), .ZN(sub_332_carry[1]) );
  INVD1 U3172 ( .I(xi4_r[48]), .ZN(n1191) );
  INVD1 U3173 ( .I(xi4_r[49]), .ZN(n1190) );
  INVD1 U3174 ( .I(xi4_r[50]), .ZN(n1189) );
  INVD1 U3175 ( .I(xi4_r[51]), .ZN(n1188) );
  INVD1 U3176 ( .I(xi4_r[52]), .ZN(n1187) );
  INVD1 U3177 ( .I(xi4_r[53]), .ZN(n1186) );
  INVD1 U3178 ( .I(xi4_r[54]), .ZN(n1185) );
  INVD1 U3179 ( .I(xi4_r[55]), .ZN(n1184) );
  INVD1 U3180 ( .I(xi4_r[56]), .ZN(n1183) );
  INVD1 U3181 ( .I(xi4_r[57]), .ZN(n1182) );
  INVD1 U3182 ( .I(xi4_r[58]), .ZN(n1181) );
  INVD1 U3183 ( .I(xi4_r[59]), .ZN(n1180) );
  INVD1 U3184 ( .I(xi4_r[60]), .ZN(n1179) );
  INVD1 U3185 ( .I(xi4_r[61]), .ZN(n1178) );
  INVD1 U3186 ( .I(xi4_r[62]), .ZN(n1177) );
  INVD1 U3187 ( .I(xi6_r[63]), .ZN(n1208) );
  OA22D0 U3188 ( .A1(n2308), .A2(n2307), .B1(n2306), .B2(n2305), .Z(n2315) );
  OA22D0 U3189 ( .A1(n2156), .A2(n2155), .B1(n2154), .B2(n2153), .Z(n2163) );
  OA22D0 U3190 ( .A1(n1982), .A2(n1981), .B1(n1980), .B2(n1979), .Z(n1989) );
  OA22D0 U3191 ( .A1(n2959), .A2(n2958), .B1(n2957), .B2(n2956), .Z(n2966) );
  OA22D0 U3192 ( .A1(n2807), .A2(n2806), .B1(n2805), .B2(n2804), .Z(n2814) );
  OA22D0 U3193 ( .A1(n2633), .A2(n2632), .B1(n2631), .B2(n2630), .Z(n2640) );
  INVD1 U3194 ( .I(xi6_i[63]), .ZN(n1338) );
  INVD1 U3195 ( .I(xi4_i[63]), .ZN(n1306) );
  INVD1 U3196 ( .I(xi4_r[63]), .ZN(n1176) );
  INVD1 U3197 ( .I(xo2_i_w_d1r[0]), .ZN(n1541) );
  INVD1 U3198 ( .I(xo2_r_w_d1r[0]), .ZN(n1525) );
  INVD1 U3199 ( .I(xo6_r_w_d1r[0]), .ZN(n1653) );
  INVD1 U3200 ( .I(xo6_i_w_d1r[0]), .ZN(n1669) );
  INVD1 U3201 ( .I(xo3_i_w_d1r[0]), .ZN(n1557) );
  INVD1 U3202 ( .I(xo7_i_w_d1r[0]), .ZN(n1685) );
  INVD1 U3203 ( .I(xo1_r_w_d1r[0]), .ZN(n1477) );
  INVD1 U3204 ( .I(xo5_r_w_d1r[0]), .ZN(n1605) );
  INVD1 U3205 ( .I(W3_8_r[55]), .ZN(n1392) );
  INVD1 U3206 ( .I(W3_8_r[54]), .ZN(n1393) );
  INVD1 U3207 ( .I(W1_8_r[55]), .ZN(n1377) );
  INVD1 U3208 ( .I(W1_8_r[54]), .ZN(n1378) );
  INVD1 U3209 ( .I(W3_8_i[56]), .ZN(n1421) );
  INVD1 U3210 ( .I(W3_8_r[56]), .ZN(n1391) );
  INVD1 U3211 ( .I(W1_8_i[56]), .ZN(n1406) );
  INVD1 U3212 ( .I(W1_8_r[56]), .ZN(n1376) );
  INVD1 U3213 ( .I(W3_8_i[57]), .ZN(n1420) );
  INVD1 U3214 ( .I(W3_8_r[57]), .ZN(n1390) );
  INVD1 U3215 ( .I(W1_8_i[57]), .ZN(n1405) );
  INVD1 U3216 ( .I(W1_8_r[57]), .ZN(n1375) );
  INVD1 U3217 ( .I(W3_8_i[58]), .ZN(n1419) );
  INVD1 U3218 ( .I(W3_8_r[58]), .ZN(n1389) );
  INVD1 U3219 ( .I(W1_8_i[58]), .ZN(n1404) );
  INVD1 U3220 ( .I(W1_8_r[58]), .ZN(n1374) );
  INVD1 U3221 ( .I(W3_8_i[59]), .ZN(n1418) );
  INVD1 U3222 ( .I(W3_8_r[59]), .ZN(n1388) );
  INVD1 U3223 ( .I(W1_8_i[59]), .ZN(n1403) );
  INVD1 U3224 ( .I(W1_8_r[59]), .ZN(n1373) );
  INVD1 U3225 ( .I(W3_8_r[49]), .ZN(n1398) );
  INVD1 U3226 ( .I(W1_8_r[49]), .ZN(n1383) );
  INVD1 U3227 ( .I(W3_8_i[49]), .ZN(n1428) );
  INVD1 U3228 ( .I(W3_8_r[50]), .ZN(n1397) );
  INVD1 U3229 ( .I(W1_8_i[49]), .ZN(n1413) );
  INVD1 U3230 ( .I(W1_8_r[50]), .ZN(n1382) );
  INVD1 U3231 ( .I(W3_8_i[50]), .ZN(n1427) );
  INVD1 U3232 ( .I(W1_8_i[50]), .ZN(n1412) );
  INVD1 U3233 ( .I(W3_8_r[51]), .ZN(n1396) );
  INVD1 U3234 ( .I(W3_8_r[52]), .ZN(n1395) );
  INVD1 U3235 ( .I(W1_8_r[51]), .ZN(n1381) );
  INVD1 U3236 ( .I(W1_8_r[52]), .ZN(n1380) );
  INVD1 U3237 ( .I(W3_8_r[53]), .ZN(n1394) );
  INVD1 U3238 ( .I(W1_8_r[53]), .ZN(n1379) );
  INVD1 U3239 ( .I(W3_8_i[51]), .ZN(n1426) );
  INVD1 U3240 ( .I(W1_8_i[51]), .ZN(n1411) );
  INVD1 U3241 ( .I(W3_8_i[52]), .ZN(n1425) );
  INVD1 U3242 ( .I(W3_8_i[53]), .ZN(n1424) );
  INVD1 U3243 ( .I(W1_8_i[52]), .ZN(n1410) );
  INVD1 U3244 ( .I(W1_8_i[53]), .ZN(n1409) );
  INVD1 U3245 ( .I(W3_8_i[55]), .ZN(n1422) );
  INVD1 U3246 ( .I(W3_8_i[54]), .ZN(n1423) );
  INVD1 U3247 ( .I(W1_8_i[55]), .ZN(n1407) );
  INVD1 U3248 ( .I(W1_8_i[54]), .ZN(n1408) );
  INVD1 U3249 ( .I(W3_8_i[60]), .ZN(n1417) );
  INVD1 U3250 ( .I(W3_8_r[60]), .ZN(n1387) );
  INVD1 U3251 ( .I(W1_8_i[60]), .ZN(n1402) );
  INVD1 U3252 ( .I(W1_8_r[60]), .ZN(n1372) );
  INVD1 U3253 ( .I(W3_8_i[61]), .ZN(n1416) );
  INVD1 U3254 ( .I(W3_8_r[61]), .ZN(n1386) );
  INVD1 U3255 ( .I(W1_8_i[61]), .ZN(n1401) );
  INVD1 U3256 ( .I(W1_8_r[61]), .ZN(n1371) );
  INVD1 U3257 ( .I(W3_8_i[62]), .ZN(n1415) );
  INVD1 U3258 ( .I(W3_8_r[62]), .ZN(n1385) );
  INVD1 U3259 ( .I(W1_8_i[62]), .ZN(n1400) );
  INVD1 U3260 ( .I(W1_8_r[62]), .ZN(n1370) );
  TIEL U3261 ( .ZN(xo7_i[0]) );
  XNR2D1 U3262 ( .A1(n1477), .A2(xo3_r_w_d1r[0]), .ZN(s2_3_tmp_i_0_) );
  XNR2D1 U3263 ( .A1(n1605), .A2(xo7_r_w_d1r[0]), .ZN(s2_7_tmp_i_0_) );
  XNR2D1 U3264 ( .A1(n1604), .A2(s2_6_i[0]), .ZN(s3_7_i[0]) );
  XNR2D1 U3265 ( .A1(n1636), .A2(s2_4_i[0]), .ZN(s3_5_i[0]) );
  XNR2D1 U3266 ( .A1(n1476), .A2(s2_2_i[0]), .ZN(s3_3_i[0]) );
  XNR2D1 U3267 ( .A1(n1508), .A2(s2_0_i[0]), .ZN(s3_1_i[0]) );
  XNR2D1 U3268 ( .A1(n1637), .A2(s2_6_r[0]), .ZN(s3_7_r[0]) );
  XNR2D1 U3269 ( .A1(n1603), .A2(s2_4_r[0]), .ZN(s3_5_r[0]) );
  XNR2D1 U3270 ( .A1(n1509), .A2(s2_2_r[0]), .ZN(s3_3_r[0]) );
  XNR2D1 U3271 ( .A1(n1475), .A2(s2_0_r[0]), .ZN(s3_1_r[0]) );
  XNR2D1 U3272 ( .A1(n1685), .A2(xo5_i_w_d1r[0]), .ZN(s2_7_i[0]) );
  XNR2D1 U3273 ( .A1(n1669), .A2(xo4_i_w_d1r[0]), .ZN(s2_6_i[0]) );
  XNR2D1 U3274 ( .A1(n1557), .A2(xo1_i_w_d1r[0]), .ZN(s2_3_i[0]) );
  XNR2D1 U3275 ( .A1(n1541), .A2(xo0_i_w_d1r[0]), .ZN(s2_2_i[0]) );
  XNR2D1 U3276 ( .A1(n1653), .A2(xo4_r_w_d1r[0]), .ZN(s2_6_r[0]) );
  XNR2D1 U3277 ( .A1(n1525), .A2(xo0_r_w_d1r[0]), .ZN(s2_2_r[0]) );
  CKXOR2D1 U3278 ( .A1(n1151), .A2(n1150), .Z(s1_6_tmp_i[1]) );
  CKXOR2D1 U3279 ( .A1(n935), .A2(n1149), .Z(s1_6_tmp_i[2]) );
  CKXOR2D1 U3280 ( .A1(n934), .A2(n1148), .Z(s1_6_tmp_i[3]) );
  CKXOR2D1 U3281 ( .A1(n923), .A2(n1147), .Z(s1_6_tmp_i[4]) );
  CKXOR2D1 U3282 ( .A1(n924), .A2(n1146), .Z(s1_6_tmp_i[5]) );
  CKXOR2D1 U3283 ( .A1(n925), .A2(n1145), .Z(s1_6_tmp_i[6]) );
  CKXOR2D1 U3284 ( .A1(n926), .A2(n1144), .Z(s1_6_tmp_i[7]) );
  CKXOR2D1 U3285 ( .A1(n927), .A2(n1143), .Z(s1_6_tmp_i[8]) );
  CKXOR2D1 U3286 ( .A1(n928), .A2(n1142), .Z(s1_6_tmp_i[9]) );
  CKXOR2D1 U3287 ( .A1(n929), .A2(n1141), .Z(s1_6_tmp_i[10]) );
  CKXOR2D1 U3288 ( .A1(n930), .A2(n1140), .Z(s1_6_tmp_i[11]) );
  CKXOR2D1 U3289 ( .A1(n931), .A2(n1139), .Z(s1_6_tmp_i[12]) );
  CKXOR2D1 U3290 ( .A1(n932), .A2(n1138), .Z(s1_6_tmp_i[13]) );
  CKXOR2D1 U3291 ( .A1(n933), .A2(n1137), .Z(s1_6_tmp_i[14]) );
  CKXOR2D1 U3292 ( .A1(s2_7_tmp_i_0_), .A2(s2_6_i[0]), .Z(s3_6_i[0]) );
  CKXOR2D1 U3293 ( .A1(s2_5_i[0]), .A2(s2_4_i[0]), .Z(s3_4_i[0]) );
  CKXOR2D1 U3294 ( .A1(s2_3_tmp_i_0_), .A2(s2_2_i[0]), .Z(s3_2_i[0]) );
  CKXOR2D1 U3295 ( .A1(s2_1_i[0]), .A2(s2_0_i[0]), .Z(s3_0_i[0]) );
  CKXOR2D1 U3296 ( .A1(s2_7_i[0]), .A2(s2_6_r[0]), .Z(s3_6_r[0]) );
  CKXOR2D1 U3297 ( .A1(s2_5_r[0]), .A2(s2_4_r[0]), .Z(s3_4_r[0]) );
  CKXOR2D1 U3298 ( .A1(s2_3_i[0]), .A2(s2_2_r[0]), .Z(s3_2_r[0]) );
  CKXOR2D1 U3299 ( .A1(s2_1_r[0]), .A2(s2_0_r[0]), .Z(s3_0_r[0]) );
  CKXOR2D1 U3300 ( .A1(xo7_i_w_d1r[0]), .A2(xo5_i_w_d1r[0]), .Z(s2_5_i[0]) );
  CKXOR2D1 U3301 ( .A1(xo6_i_w_d1r[0]), .A2(xo4_i_w_d1r[0]), .Z(s2_4_i[0]) );
  CKXOR2D1 U3302 ( .A1(xo3_i_w_d1r[0]), .A2(xo1_i_w_d1r[0]), .Z(s2_1_i[0]) );
  CKXOR2D1 U3303 ( .A1(xo2_i_w_d1r[0]), .A2(xo0_i_w_d1r[0]), .Z(s2_0_i[0]) );
  CKXOR2D1 U3304 ( .A1(xo7_r_w_d1r[0]), .A2(xo5_r_w_d1r[0]), .Z(s2_5_r[0]) );
  CKXOR2D1 U3305 ( .A1(xo6_r_w_d1r[0]), .A2(xo4_r_w_d1r[0]), .Z(s2_4_r[0]) );
  CKXOR2D1 U3306 ( .A1(xo3_r_w_d1r[0]), .A2(xo1_r_w_d1r[0]), .Z(s2_1_r[0]) );
  CKXOR2D1 U3307 ( .A1(xo2_r_w_d1r[0]), .A2(xo0_r_w_d1r[0]), .Z(s2_0_r[0]) );
  AN2XD1 U3308 ( .A1(xi4_r[47]), .A2(xi0_r[47]), .Z(add_328_carry[1]) );
  AN2XD1 U3309 ( .A1(xi5_r[47]), .A2(xi1_r[47]), .Z(add_329_carry[1]) );
  AN2XD1 U3310 ( .A1(xi6_r[47]), .A2(xi2_r[47]), .Z(add_330_carry[1]) );
  AN2XD1 U3311 ( .A1(xi7_r[47]), .A2(xi3_r[47]), .Z(add_331_carry[1]) );
  AN2XD1 U3312 ( .A1(xi4_i[47]), .A2(xi0_i[47]), .Z(add_337_carry[1]) );
  AN2XD1 U3313 ( .A1(xi5_i[47]), .A2(xi1_i[47]), .Z(add_338_carry[1]) );
  AN2XD1 U3314 ( .A1(xi6_i[47]), .A2(xi2_i[47]), .Z(add_339_carry[1]) );
  AN2XD1 U3315 ( .A1(xi7_i[47]), .A2(xi3_i[47]), .Z(add_340_carry[1]) );
  XNR2D1 U3316 ( .A1(n1072), .A2(n1419), .ZN(n1724) );
  XNR2D1 U3317 ( .A1(n1073), .A2(s1_7_i[11]), .ZN(n1686) );
  XNR2D1 U3318 ( .A1(n1073), .A2(n1418), .ZN(n1723) );
  XNR2D1 U3319 ( .A1(s1_7_i[6]), .A2(W3_8_i[63]), .ZN(n1767) );
  XNR2D1 U3320 ( .A1(n1080), .A2(n1415), .ZN(n1768) );
  XNR2D1 U3321 ( .A1(n1081), .A2(s1_7_i[5]), .ZN(n1687) );
  XNR2D1 U3322 ( .A1(s1_7_i[4]), .A2(W3_8_i[63]), .ZN(n1785) );
  XNR2D1 U3323 ( .A1(n1084), .A2(n1415), .ZN(n1786) );
  XNR2D1 U3324 ( .A1(n1085), .A2(s1_7_i[3]), .ZN(n1688) );
  XNR2D1 U3325 ( .A1(n1077), .A2(n1420), .ZN(n1755) );
  XNR2D1 U3326 ( .A1(n1078), .A2(s1_7_i[7]), .ZN(n1689) );
  XNR2D1 U3327 ( .A1(n1079), .A2(n1419), .ZN(n1754) );
  XNR2D1 U3328 ( .A1(n1069), .A2(n1426), .ZN(n1717) );
  XNR2D1 U3329 ( .A1(n1070), .A2(s1_7_i[13]), .ZN(n1690) );
  XNR2D1 U3330 ( .A1(n1071), .A2(n1425), .ZN(n1716) );
  XNR2D1 U3331 ( .A1(n1692), .A2(n1691), .ZN(dp_cluster_0_mult_486_C412_n162)
         );
  XNR2D1 U3332 ( .A1(n1067), .A2(s1_7_i[15]), .ZN(n1693) );
  XNR2D1 U3333 ( .A1(n1075), .A2(s1_7_i[9]), .ZN(n1694) );
  XNR2D1 U3334 ( .A1(n1068), .A2(n1418), .ZN(n1695) );
  XNR2D1 U3335 ( .A1(s1_7_i[16]), .A2(W3_8_i[60]), .ZN(n1827) );
  XNR2D1 U3336 ( .A1(n1068), .A2(n1419), .ZN(n1696) );
  XNR2D1 U3337 ( .A1(n1068), .A2(n1420), .ZN(n1697) );
  XNR2D1 U3338 ( .A1(n1068), .A2(n1421), .ZN(n1698) );
  XNR2D1 U3339 ( .A1(n1068), .A2(n1422), .ZN(n1699) );
  XNR2D1 U3340 ( .A1(n1068), .A2(n1423), .ZN(n1700) );
  XNR2D1 U3341 ( .A1(n1068), .A2(n1424), .ZN(n1701) );
  XNR2D1 U3342 ( .A1(n1068), .A2(n1425), .ZN(n1702) );
  XNR2D1 U3343 ( .A1(n1068), .A2(n1426), .ZN(n1703) );
  XNR2D1 U3344 ( .A1(n1068), .A2(n1427), .ZN(n1704) );
  XNR2D1 U3345 ( .A1(n1068), .A2(n1428), .ZN(n1705) );
  XNR2D1 U3346 ( .A1(n1100), .A2(n1068), .ZN(n1706) );
  XNR2D1 U3347 ( .A1(n1070), .A2(n1416), .ZN(n1707) );
  XNR2D1 U3348 ( .A1(n1070), .A2(n1415), .ZN(n1834) );
  XNR2D1 U3349 ( .A1(n1070), .A2(n1417), .ZN(n1708) );
  XNR2D1 U3350 ( .A1(n1070), .A2(n1418), .ZN(n1709) );
  XNR2D1 U3351 ( .A1(n1070), .A2(n1419), .ZN(n1710) );
  XNR2D1 U3352 ( .A1(n1070), .A2(n1420), .ZN(n1711) );
  XNR2D1 U3353 ( .A1(n1070), .A2(n1421), .ZN(n1712) );
  XNR2D1 U3354 ( .A1(n1070), .A2(n1422), .ZN(n1713) );
  XNR2D1 U3355 ( .A1(n1070), .A2(n1423), .ZN(n1714) );
  XNR2D1 U3356 ( .A1(n1070), .A2(n1424), .ZN(n1715) );
  XNR2D1 U3357 ( .A1(n1070), .A2(n1427), .ZN(n1718) );
  XNR2D1 U3358 ( .A1(n1070), .A2(n1428), .ZN(n1719) );
  XNR2D1 U3359 ( .A1(n1100), .A2(n1071), .ZN(n1720) );
  XNR2D1 U3360 ( .A1(s1_7_i[12]), .A2(W3_8_i[63]), .ZN(n1821) );
  AO21D1 U3361 ( .A1(n953), .A2(n1822), .B(n1821), .Z(
        dp_cluster_0_mult_486_C412_n281) );
  XNR2D1 U3362 ( .A1(n1073), .A2(n1416), .ZN(n1721) );
  XNR2D1 U3363 ( .A1(n1073), .A2(n1415), .ZN(n1820) );
  XNR2D1 U3364 ( .A1(n1073), .A2(n1417), .ZN(n1722) );
  XNR2D1 U3365 ( .A1(n1073), .A2(n1420), .ZN(n1725) );
  XNR2D1 U3366 ( .A1(n1073), .A2(n1421), .ZN(n1726) );
  XNR2D1 U3367 ( .A1(n1073), .A2(n1422), .ZN(n1727) );
  XNR2D1 U3368 ( .A1(n1073), .A2(n1423), .ZN(n1728) );
  XNR2D1 U3369 ( .A1(n1073), .A2(n1424), .ZN(n1729) );
  XNR2D1 U3370 ( .A1(n1073), .A2(n1425), .ZN(n1730) );
  XNR2D1 U3371 ( .A1(n1073), .A2(n1426), .ZN(n1731) );
  XNR2D1 U3372 ( .A1(n1073), .A2(n1427), .ZN(n1732) );
  XNR2D1 U3373 ( .A1(n1073), .A2(n1428), .ZN(n1733) );
  XNR2D1 U3374 ( .A1(n1100), .A2(n1073), .ZN(n1734) );
  XNR2D1 U3375 ( .A1(s1_7_i[10]), .A2(W3_8_i[63]), .ZN(n1825) );
  AO21D1 U3376 ( .A1(n958), .A2(n1826), .B(n1825), .Z(
        dp_cluster_0_mult_486_C412_n296) );
  XNR2D1 U3377 ( .A1(n1076), .A2(n1416), .ZN(n1735) );
  XNR2D1 U3378 ( .A1(n1075), .A2(n1415), .ZN(n1824) );
  XNR2D1 U3379 ( .A1(n1075), .A2(n1417), .ZN(n1736) );
  XNR2D1 U3380 ( .A1(n1075), .A2(n1418), .ZN(n1737) );
  XNR2D1 U3381 ( .A1(n1075), .A2(n1419), .ZN(n1738) );
  XNR2D1 U3382 ( .A1(n1075), .A2(n1420), .ZN(n1739) );
  XNR2D1 U3383 ( .A1(n1075), .A2(n1421), .ZN(n1740) );
  XNR2D1 U3384 ( .A1(n1075), .A2(n1422), .ZN(n1741) );
  XNR2D1 U3385 ( .A1(n1075), .A2(n1423), .ZN(n1742) );
  XNR2D1 U3386 ( .A1(n1075), .A2(n1424), .ZN(n1743) );
  XNR2D1 U3387 ( .A1(n1075), .A2(n1425), .ZN(n1744) );
  XNR2D1 U3388 ( .A1(n1075), .A2(n1426), .ZN(n1745) );
  XNR2D1 U3389 ( .A1(n1075), .A2(n1427), .ZN(n1746) );
  XNR2D1 U3390 ( .A1(n1075), .A2(n1428), .ZN(n1747) );
  XNR2D1 U3391 ( .A1(n1100), .A2(n1076), .ZN(n1748) );
  XNR2D1 U3392 ( .A1(s1_7_i[8]), .A2(W3_8_i[63]), .ZN(n1749) );
  AO21D1 U3393 ( .A1(n956), .A2(n1766), .B(n1749), .Z(
        dp_cluster_0_mult_486_C412_n312) );
  XNR2D1 U3394 ( .A1(n1078), .A2(n1415), .ZN(n1750) );
  XNR2D1 U3395 ( .A1(n1078), .A2(n1416), .ZN(n1751) );
  XNR2D1 U3396 ( .A1(n1078), .A2(n1417), .ZN(n1752) );
  XNR2D1 U3397 ( .A1(n1078), .A2(n1418), .ZN(n1753) );
  XNR2D1 U3398 ( .A1(n1078), .A2(n1421), .ZN(n1756) );
  XNR2D1 U3399 ( .A1(n1078), .A2(n1422), .ZN(n1757) );
  XNR2D1 U3400 ( .A1(n1078), .A2(n1423), .ZN(n1758) );
  XNR2D1 U3401 ( .A1(n1078), .A2(n1424), .ZN(n1759) );
  XNR2D1 U3402 ( .A1(n1078), .A2(n1425), .ZN(n1760) );
  XNR2D1 U3403 ( .A1(n1078), .A2(n1426), .ZN(n1761) );
  XNR2D1 U3404 ( .A1(n1078), .A2(n1427), .ZN(n1762) );
  XNR2D1 U3405 ( .A1(n1078), .A2(n1428), .ZN(n1763) );
  XNR2D1 U3406 ( .A1(n1099), .A2(n1079), .ZN(n1765) );
  AO21D1 U3407 ( .A1(n954), .A2(n1784), .B(n1767), .Z(
        dp_cluster_0_mult_486_C412_n329) );
  XNR2D1 U3408 ( .A1(n1081), .A2(n1416), .ZN(n1769) );
  XNR2D1 U3409 ( .A1(n1081), .A2(n1417), .ZN(n1770) );
  XNR2D1 U3410 ( .A1(n1081), .A2(n1418), .ZN(n1771) );
  XNR2D1 U3411 ( .A1(n1081), .A2(n1419), .ZN(n1772) );
  XNR2D1 U3412 ( .A1(n1081), .A2(n1420), .ZN(n1773) );
  XNR2D1 U3413 ( .A1(n1081), .A2(n1421), .ZN(n1774) );
  XNR2D1 U3414 ( .A1(n1081), .A2(n1422), .ZN(n1775) );
  XNR2D1 U3415 ( .A1(n1081), .A2(n1423), .ZN(n1776) );
  XNR2D1 U3416 ( .A1(n1081), .A2(n1424), .ZN(n1777) );
  XNR2D1 U3417 ( .A1(n1081), .A2(n1425), .ZN(n1778) );
  XNR2D1 U3418 ( .A1(n1081), .A2(n1426), .ZN(n1779) );
  XNR2D1 U3419 ( .A1(n1081), .A2(n1427), .ZN(n1780) );
  XNR2D1 U3420 ( .A1(n1081), .A2(n1428), .ZN(n1781) );
  XNR2D1 U3421 ( .A1(n1099), .A2(n1082), .ZN(n1783) );
  AO21D1 U3422 ( .A1(n955), .A2(n1802), .B(n1785), .Z(
        dp_cluster_0_mult_486_C412_n345) );
  XNR2D1 U3423 ( .A1(n1084), .A2(n1416), .ZN(n1787) );
  XNR2D1 U3424 ( .A1(n1084), .A2(n1417), .ZN(n1788) );
  XNR2D1 U3425 ( .A1(n1084), .A2(n1418), .ZN(n1789) );
  XNR2D1 U3426 ( .A1(n1084), .A2(n1419), .ZN(n1790) );
  XNR2D1 U3427 ( .A1(n1084), .A2(n1420), .ZN(n1791) );
  XNR2D1 U3428 ( .A1(n1084), .A2(n1421), .ZN(n1792) );
  XNR2D1 U3429 ( .A1(n1084), .A2(n1422), .ZN(n1793) );
  XNR2D1 U3430 ( .A1(n1084), .A2(n1423), .ZN(n1794) );
  XNR2D1 U3431 ( .A1(n1084), .A2(n1424), .ZN(n1795) );
  XNR2D1 U3432 ( .A1(n1084), .A2(n1425), .ZN(n1796) );
  XNR2D1 U3433 ( .A1(n1084), .A2(n1426), .ZN(n1797) );
  XNR2D1 U3434 ( .A1(n1084), .A2(n1427), .ZN(n1798) );
  XNR2D1 U3435 ( .A1(n1084), .A2(n1428), .ZN(n1799) );
  XNR2D1 U3436 ( .A1(n1099), .A2(n1085), .ZN(n1801) );
  CKXOR2D1 U3437 ( .A1(n1103), .A2(W3_8_i[63]), .Z(n1803) );
  XNR2D1 U3438 ( .A1(n1103), .A2(W3_8_i[62]), .ZN(n1804) );
  MOAI22D1 U3439 ( .A1(n1804), .A2(n1818), .B1(n1803), .B2(s1_7_i[1]), .ZN(
        dp_cluster_0_mult_486_C412_n362) );
  XNR2D1 U3440 ( .A1(n1102), .A2(W3_8_i[61]), .ZN(n1805) );
  XNR2D1 U3441 ( .A1(n1103), .A2(W3_8_i[60]), .ZN(n1806) );
  XNR2D1 U3442 ( .A1(n1103), .A2(W3_8_i[59]), .ZN(n1807) );
  XNR2D1 U3443 ( .A1(n1102), .A2(W3_8_i[58]), .ZN(n1808) );
  XNR2D1 U3444 ( .A1(n1102), .A2(W3_8_i[57]), .ZN(n1809) );
  XNR2D1 U3445 ( .A1(n1102), .A2(W3_8_i[56]), .ZN(n1810) );
  XNR2D1 U3446 ( .A1(n1102), .A2(W3_8_i[55]), .ZN(n1811) );
  XNR2D1 U3447 ( .A1(n1102), .A2(W3_8_i[54]), .ZN(n1812) );
  XNR2D1 U3448 ( .A1(n1102), .A2(W3_8_i[53]), .ZN(n1813) );
  XNR2D1 U3449 ( .A1(n1102), .A2(W3_8_i[52]), .ZN(n1814) );
  XNR2D1 U3450 ( .A1(n1102), .A2(W3_8_i[51]), .ZN(n1815) );
  XNR2D1 U3451 ( .A1(n1102), .A2(W3_8_i[50]), .ZN(n1816) );
  XNR2D1 U3452 ( .A1(n1102), .A2(W3_8_i[49]), .ZN(n1817) );
  XNR2D1 U3453 ( .A1(W3_8_i[61]), .A2(s1_7_i[16]), .ZN(n1830) );
  XNR2D1 U3454 ( .A1(s1_7_i[14]), .A2(W3_8_i[63]), .ZN(n1831) );
  XNR2D1 U3455 ( .A1(n1028), .A2(n1389), .ZN(n1876) );
  XNR2D1 U3456 ( .A1(n1029), .A2(s1_7_r[11]), .ZN(n1838) );
  XNR2D1 U3457 ( .A1(n1029), .A2(n1388), .ZN(n1875) );
  XNR2D1 U3458 ( .A1(s1_7_r[6]), .A2(W3_8_r[63]), .ZN(n1919) );
  XNR2D1 U3459 ( .A1(n1036), .A2(n1385), .ZN(n1920) );
  XNR2D1 U3460 ( .A1(n1037), .A2(s1_7_r[5]), .ZN(n1839) );
  XNR2D1 U3461 ( .A1(s1_7_r[4]), .A2(W3_8_r[63]), .ZN(n1937) );
  XNR2D1 U3462 ( .A1(n1040), .A2(n1385), .ZN(n1938) );
  XNR2D1 U3463 ( .A1(n1041), .A2(s1_7_r[3]), .ZN(n1840) );
  XNR2D1 U3464 ( .A1(n1033), .A2(n1390), .ZN(n1907) );
  XNR2D1 U3465 ( .A1(n1034), .A2(s1_7_r[7]), .ZN(n1841) );
  XNR2D1 U3466 ( .A1(n1035), .A2(n1389), .ZN(n1906) );
  XNR2D1 U3467 ( .A1(n1025), .A2(n1396), .ZN(n1869) );
  XNR2D1 U3468 ( .A1(n1026), .A2(s1_7_r[13]), .ZN(n1842) );
  XNR2D1 U3469 ( .A1(n1027), .A2(n1395), .ZN(n1868) );
  XNR2D1 U3470 ( .A1(n1844), .A2(n1843), .ZN(dp_cluster_0_mult_485_C412_n162)
         );
  XNR2D1 U3471 ( .A1(n1023), .A2(s1_7_r[15]), .ZN(n1845) );
  XNR2D1 U3472 ( .A1(n1031), .A2(s1_7_r[9]), .ZN(n1846) );
  XNR2D1 U3473 ( .A1(n1024), .A2(n1388), .ZN(n1847) );
  XNR2D1 U3474 ( .A1(s1_7_r[16]), .A2(W3_8_r[60]), .ZN(n1979) );
  XNR2D1 U3475 ( .A1(n1024), .A2(n1389), .ZN(n1848) );
  XNR2D1 U3476 ( .A1(n1024), .A2(n1390), .ZN(n1849) );
  XNR2D1 U3477 ( .A1(n1024), .A2(n1391), .ZN(n1850) );
  XNR2D1 U3478 ( .A1(n1024), .A2(n1392), .ZN(n1851) );
  XNR2D1 U3479 ( .A1(n1024), .A2(n1393), .ZN(n1852) );
  XNR2D1 U3480 ( .A1(n1024), .A2(n1394), .ZN(n1853) );
  XNR2D1 U3481 ( .A1(n1024), .A2(n1395), .ZN(n1854) );
  XNR2D1 U3482 ( .A1(n1024), .A2(n1396), .ZN(n1855) );
  XNR2D1 U3483 ( .A1(n1024), .A2(n1397), .ZN(n1856) );
  XNR2D1 U3484 ( .A1(n1024), .A2(n1398), .ZN(n1857) );
  XNR2D1 U3485 ( .A1(n1094), .A2(n1024), .ZN(n1858) );
  XNR2D1 U3486 ( .A1(n1026), .A2(n1386), .ZN(n1859) );
  XNR2D1 U3487 ( .A1(n1026), .A2(n1385), .ZN(n1986) );
  XNR2D1 U3488 ( .A1(n1026), .A2(n1387), .ZN(n1860) );
  XNR2D1 U3489 ( .A1(n1026), .A2(n1388), .ZN(n1861) );
  XNR2D1 U3490 ( .A1(n1026), .A2(n1389), .ZN(n1862) );
  XNR2D1 U3491 ( .A1(n1026), .A2(n1390), .ZN(n1863) );
  XNR2D1 U3492 ( .A1(n1026), .A2(n1391), .ZN(n1864) );
  XNR2D1 U3493 ( .A1(n1026), .A2(n1392), .ZN(n1865) );
  XNR2D1 U3494 ( .A1(n1026), .A2(n1393), .ZN(n1866) );
  XNR2D1 U3495 ( .A1(n1026), .A2(n1394), .ZN(n1867) );
  XNR2D1 U3496 ( .A1(n1026), .A2(n1397), .ZN(n1870) );
  XNR2D1 U3497 ( .A1(n1026), .A2(n1398), .ZN(n1871) );
  XNR2D1 U3498 ( .A1(n1094), .A2(n1027), .ZN(n1872) );
  XNR2D1 U3499 ( .A1(s1_7_r[12]), .A2(W3_8_r[63]), .ZN(n1973) );
  AO21D1 U3500 ( .A1(n959), .A2(n1974), .B(n1973), .Z(
        dp_cluster_0_mult_485_C412_n281) );
  XNR2D1 U3501 ( .A1(n1029), .A2(n1386), .ZN(n1873) );
  XNR2D1 U3502 ( .A1(n1029), .A2(n1385), .ZN(n1972) );
  XNR2D1 U3503 ( .A1(n1029), .A2(n1387), .ZN(n1874) );
  XNR2D1 U3504 ( .A1(n1029), .A2(n1390), .ZN(n1877) );
  XNR2D1 U3505 ( .A1(n1029), .A2(n1391), .ZN(n1878) );
  XNR2D1 U3506 ( .A1(n1029), .A2(n1392), .ZN(n1879) );
  XNR2D1 U3507 ( .A1(n1029), .A2(n1393), .ZN(n1880) );
  XNR2D1 U3508 ( .A1(n1029), .A2(n1394), .ZN(n1881) );
  XNR2D1 U3509 ( .A1(n1029), .A2(n1395), .ZN(n1882) );
  XNR2D1 U3510 ( .A1(n1029), .A2(n1396), .ZN(n1883) );
  XNR2D1 U3511 ( .A1(n1029), .A2(n1397), .ZN(n1884) );
  XNR2D1 U3512 ( .A1(n1029), .A2(n1398), .ZN(n1885) );
  XNR2D1 U3513 ( .A1(n1094), .A2(n1029), .ZN(n1886) );
  XNR2D1 U3514 ( .A1(s1_7_r[10]), .A2(W3_8_r[63]), .ZN(n1977) );
  AO21D1 U3515 ( .A1(n964), .A2(n1978), .B(n1977), .Z(
        dp_cluster_0_mult_485_C412_n296) );
  XNR2D1 U3516 ( .A1(n1032), .A2(n1386), .ZN(n1887) );
  XNR2D1 U3517 ( .A1(n1031), .A2(n1385), .ZN(n1976) );
  XNR2D1 U3518 ( .A1(n1031), .A2(n1387), .ZN(n1888) );
  XNR2D1 U3519 ( .A1(n1031), .A2(n1388), .ZN(n1889) );
  XNR2D1 U3520 ( .A1(n1031), .A2(n1389), .ZN(n1890) );
  XNR2D1 U3521 ( .A1(n1031), .A2(n1390), .ZN(n1891) );
  XNR2D1 U3522 ( .A1(n1031), .A2(n1391), .ZN(n1892) );
  XNR2D1 U3523 ( .A1(n1031), .A2(n1392), .ZN(n1893) );
  XNR2D1 U3524 ( .A1(n1031), .A2(n1393), .ZN(n1894) );
  XNR2D1 U3525 ( .A1(n1031), .A2(n1394), .ZN(n1895) );
  XNR2D1 U3526 ( .A1(n1031), .A2(n1395), .ZN(n1896) );
  XNR2D1 U3527 ( .A1(n1031), .A2(n1396), .ZN(n1897) );
  XNR2D1 U3528 ( .A1(n1031), .A2(n1397), .ZN(n1898) );
  XNR2D1 U3529 ( .A1(n1031), .A2(n1398), .ZN(n1899) );
  XNR2D1 U3530 ( .A1(n1094), .A2(n1032), .ZN(n1900) );
  XNR2D1 U3531 ( .A1(s1_7_r[8]), .A2(W3_8_r[63]), .ZN(n1901) );
  AO21D1 U3532 ( .A1(n962), .A2(n1918), .B(n1901), .Z(
        dp_cluster_0_mult_485_C412_n312) );
  XNR2D1 U3533 ( .A1(n1034), .A2(n1385), .ZN(n1902) );
  XNR2D1 U3534 ( .A1(n1034), .A2(n1386), .ZN(n1903) );
  XNR2D1 U3535 ( .A1(n1034), .A2(n1387), .ZN(n1904) );
  XNR2D1 U3536 ( .A1(n1034), .A2(n1388), .ZN(n1905) );
  XNR2D1 U3537 ( .A1(n1034), .A2(n1391), .ZN(n1908) );
  XNR2D1 U3538 ( .A1(n1034), .A2(n1392), .ZN(n1909) );
  XNR2D1 U3539 ( .A1(n1034), .A2(n1393), .ZN(n1910) );
  XNR2D1 U3540 ( .A1(n1034), .A2(n1394), .ZN(n1911) );
  XNR2D1 U3541 ( .A1(n1034), .A2(n1395), .ZN(n1912) );
  XNR2D1 U3542 ( .A1(n1034), .A2(n1396), .ZN(n1913) );
  XNR2D1 U3543 ( .A1(n1034), .A2(n1397), .ZN(n1914) );
  XNR2D1 U3544 ( .A1(n1034), .A2(n1398), .ZN(n1915) );
  XNR2D1 U3545 ( .A1(n1093), .A2(n1035), .ZN(n1917) );
  AO21D1 U3546 ( .A1(n960), .A2(n1936), .B(n1919), .Z(
        dp_cluster_0_mult_485_C412_n329) );
  XNR2D1 U3547 ( .A1(n1037), .A2(n1386), .ZN(n1921) );
  XNR2D1 U3548 ( .A1(n1037), .A2(n1387), .ZN(n1922) );
  XNR2D1 U3549 ( .A1(n1037), .A2(n1388), .ZN(n1923) );
  XNR2D1 U3550 ( .A1(n1037), .A2(n1389), .ZN(n1924) );
  XNR2D1 U3551 ( .A1(n1037), .A2(n1390), .ZN(n1925) );
  XNR2D1 U3552 ( .A1(n1037), .A2(n1391), .ZN(n1926) );
  XNR2D1 U3553 ( .A1(n1037), .A2(n1392), .ZN(n1927) );
  XNR2D1 U3554 ( .A1(n1037), .A2(n1393), .ZN(n1928) );
  XNR2D1 U3555 ( .A1(n1037), .A2(n1394), .ZN(n1929) );
  XNR2D1 U3556 ( .A1(n1037), .A2(n1395), .ZN(n1930) );
  XNR2D1 U3557 ( .A1(n1037), .A2(n1396), .ZN(n1931) );
  XNR2D1 U3558 ( .A1(n1037), .A2(n1397), .ZN(n1932) );
  XNR2D1 U3559 ( .A1(n1037), .A2(n1398), .ZN(n1933) );
  XNR2D1 U3560 ( .A1(n1093), .A2(n1038), .ZN(n1935) );
  AO21D1 U3561 ( .A1(n961), .A2(n1954), .B(n1937), .Z(
        dp_cluster_0_mult_485_C412_n345) );
  XNR2D1 U3562 ( .A1(n1040), .A2(n1386), .ZN(n1939) );
  XNR2D1 U3563 ( .A1(n1040), .A2(n1387), .ZN(n1940) );
  XNR2D1 U3564 ( .A1(n1040), .A2(n1388), .ZN(n1941) );
  XNR2D1 U3565 ( .A1(n1040), .A2(n1389), .ZN(n1942) );
  XNR2D1 U3566 ( .A1(n1040), .A2(n1390), .ZN(n1943) );
  XNR2D1 U3567 ( .A1(n1040), .A2(n1391), .ZN(n1944) );
  XNR2D1 U3568 ( .A1(n1040), .A2(n1392), .ZN(n1945) );
  XNR2D1 U3569 ( .A1(n1040), .A2(n1393), .ZN(n1946) );
  XNR2D1 U3570 ( .A1(n1040), .A2(n1394), .ZN(n1947) );
  XNR2D1 U3571 ( .A1(n1040), .A2(n1395), .ZN(n1948) );
  XNR2D1 U3572 ( .A1(n1040), .A2(n1396), .ZN(n1949) );
  XNR2D1 U3573 ( .A1(n1040), .A2(n1397), .ZN(n1950) );
  XNR2D1 U3574 ( .A1(n1040), .A2(n1398), .ZN(n1951) );
  XNR2D1 U3575 ( .A1(n1093), .A2(n1041), .ZN(n1953) );
  CKXOR2D1 U3576 ( .A1(n1109), .A2(W3_8_r[63]), .Z(n1955) );
  XNR2D1 U3577 ( .A1(n1109), .A2(W3_8_r[62]), .ZN(n1956) );
  MOAI22D1 U3578 ( .A1(n1956), .A2(n1970), .B1(n1955), .B2(s1_7_r[1]), .ZN(
        dp_cluster_0_mult_485_C412_n362) );
  XNR2D1 U3579 ( .A1(n1108), .A2(W3_8_r[61]), .ZN(n1957) );
  XNR2D1 U3580 ( .A1(n1109), .A2(W3_8_r[60]), .ZN(n1958) );
  XNR2D1 U3581 ( .A1(n1109), .A2(W3_8_r[59]), .ZN(n1959) );
  XNR2D1 U3582 ( .A1(n1108), .A2(W3_8_r[58]), .ZN(n1960) );
  XNR2D1 U3583 ( .A1(n1108), .A2(W3_8_r[57]), .ZN(n1961) );
  XNR2D1 U3584 ( .A1(n1108), .A2(W3_8_r[56]), .ZN(n1962) );
  XNR2D1 U3585 ( .A1(n1108), .A2(W3_8_r[55]), .ZN(n1963) );
  XNR2D1 U3586 ( .A1(n1108), .A2(W3_8_r[54]), .ZN(n1964) );
  XNR2D1 U3587 ( .A1(n1108), .A2(W3_8_r[53]), .ZN(n1965) );
  XNR2D1 U3588 ( .A1(n1108), .A2(W3_8_r[52]), .ZN(n1966) );
  XNR2D1 U3589 ( .A1(n1108), .A2(W3_8_r[51]), .ZN(n1967) );
  XNR2D1 U3590 ( .A1(n1108), .A2(W3_8_r[50]), .ZN(n1968) );
  XNR2D1 U3591 ( .A1(n1108), .A2(W3_8_r[49]), .ZN(n1969) );
  XNR2D1 U3592 ( .A1(W3_8_r[61]), .A2(s1_7_r[16]), .ZN(n1982) );
  XNR2D1 U3593 ( .A1(s1_7_r[14]), .A2(W3_8_r[63]), .ZN(n1983) );
  AN2XD1 U3594 ( .A1(n1991), .A2(n1174), .Z(n1990) );
  MAOI22D1 U3595 ( .A1(n1993), .A2(dp_cluster_0_N59), .B1(dp_cluster_0_N87), 
        .B2(n1992), .ZN(n1995) );
  AN2XD1 U3596 ( .A1(n1995), .A2(n1171), .Z(n1994) );
  MAOI22D1 U3597 ( .A1(n1997), .A2(dp_cluster_0_N61), .B1(dp_cluster_0_N89), 
        .B2(n1996), .ZN(n1999) );
  AN2XD1 U3598 ( .A1(n1999), .A2(n1167), .Z(n1998) );
  MAOI22D1 U3599 ( .A1(n2001), .A2(dp_cluster_0_N63), .B1(dp_cluster_0_N91), 
        .B2(n2000), .ZN(n2003) );
  AN2XD1 U3600 ( .A1(n2003), .A2(n1164), .Z(n2002) );
  MAOI22D1 U3601 ( .A1(n2005), .A2(dp_cluster_0_N65), .B1(dp_cluster_0_N93), 
        .B2(n2004), .ZN(n2007) );
  AN2XD1 U3602 ( .A1(n2007), .A2(n1160), .Z(n2006) );
  MAOI22D1 U3603 ( .A1(n2009), .A2(dp_cluster_0_N67), .B1(dp_cluster_0_N95), 
        .B2(n2008), .ZN(n2011) );
  AN2XD1 U3604 ( .A1(n2011), .A2(n1155), .Z(n2010) );
  XNR2D1 U3605 ( .A1(n1073), .A2(n1389), .ZN(n2050) );
  XNR2D1 U3606 ( .A1(n1073), .A2(s1_7_i[11]), .ZN(n2012) );
  XNR2D1 U3607 ( .A1(n1072), .A2(n1388), .ZN(n2049) );
  XNR2D1 U3608 ( .A1(s1_7_i[6]), .A2(W3_8_r[63]), .ZN(n2093) );
  XNR2D1 U3609 ( .A1(n1081), .A2(n1385), .ZN(n2094) );
  XNR2D1 U3610 ( .A1(n1081), .A2(s1_7_i[5]), .ZN(n2013) );
  XNR2D1 U3611 ( .A1(s1_7_i[4]), .A2(W3_8_r[63]), .ZN(n2111) );
  XNR2D1 U3612 ( .A1(n1084), .A2(n1385), .ZN(n2112) );
  XNR2D1 U3613 ( .A1(n1084), .A2(s1_7_i[3]), .ZN(n2014) );
  XNR2D1 U3614 ( .A1(n1078), .A2(n1390), .ZN(n2081) );
  XNR2D1 U3615 ( .A1(n1078), .A2(s1_7_i[7]), .ZN(n2015) );
  XNR2D1 U3616 ( .A1(n1078), .A2(n1389), .ZN(n2080) );
  XNR2D1 U3617 ( .A1(n1070), .A2(n1396), .ZN(n2043) );
  XNR2D1 U3618 ( .A1(n1070), .A2(s1_7_i[13]), .ZN(n2016) );
  XNR2D1 U3619 ( .A1(n1070), .A2(n1395), .ZN(n2042) );
  XNR2D1 U3620 ( .A1(n2018), .A2(n2017), .ZN(dp_cluster_1_mult_513_C418_n162)
         );
  XNR2D1 U3621 ( .A1(n1067), .A2(s1_7_i[15]), .ZN(n2019) );
  XNR2D1 U3622 ( .A1(n1075), .A2(s1_7_i[9]), .ZN(n2020) );
  XNR2D1 U3623 ( .A1(n1067), .A2(n1388), .ZN(n2021) );
  XNR2D1 U3624 ( .A1(s1_7_i[16]), .A2(W3_8_r[60]), .ZN(n2153) );
  XNR2D1 U3625 ( .A1(n1067), .A2(n1389), .ZN(n2022) );
  XNR2D1 U3626 ( .A1(n1067), .A2(n1390), .ZN(n2023) );
  XNR2D1 U3627 ( .A1(n1067), .A2(n1391), .ZN(n2024) );
  XNR2D1 U3628 ( .A1(n1067), .A2(n1392), .ZN(n2025) );
  XNR2D1 U3629 ( .A1(n1067), .A2(n1393), .ZN(n2026) );
  XNR2D1 U3630 ( .A1(n1067), .A2(n1394), .ZN(n2027) );
  XNR2D1 U3631 ( .A1(n1067), .A2(n1395), .ZN(n2028) );
  XNR2D1 U3632 ( .A1(n1067), .A2(n1396), .ZN(n2029) );
  XNR2D1 U3633 ( .A1(n1067), .A2(n1397), .ZN(n2030) );
  XNR2D1 U3634 ( .A1(n1067), .A2(n1398), .ZN(n2031) );
  XNR2D1 U3635 ( .A1(n1093), .A2(n1068), .ZN(n2032) );
  XNR2D1 U3636 ( .A1(n1069), .A2(n1386), .ZN(n2033) );
  XNR2D1 U3637 ( .A1(n1069), .A2(n1385), .ZN(n2160) );
  XNR2D1 U3638 ( .A1(n1069), .A2(n1387), .ZN(n2034) );
  XNR2D1 U3639 ( .A1(n1069), .A2(n1388), .ZN(n2035) );
  XNR2D1 U3640 ( .A1(n1070), .A2(n1389), .ZN(n2036) );
  XNR2D1 U3641 ( .A1(n1069), .A2(n1390), .ZN(n2037) );
  XNR2D1 U3642 ( .A1(n1069), .A2(n1391), .ZN(n2038) );
  XNR2D1 U3643 ( .A1(n1069), .A2(n1392), .ZN(n2039) );
  XNR2D1 U3644 ( .A1(n1069), .A2(n1393), .ZN(n2040) );
  XNR2D1 U3645 ( .A1(n1069), .A2(n1394), .ZN(n2041) );
  XNR2D1 U3646 ( .A1(n1069), .A2(n1397), .ZN(n2044) );
  XNR2D1 U3647 ( .A1(n1069), .A2(n1398), .ZN(n2045) );
  XNR2D1 U3648 ( .A1(n1092), .A2(n1071), .ZN(n2046) );
  XNR2D1 U3649 ( .A1(s1_7_i[12]), .A2(W3_8_r[63]), .ZN(n2147) );
  AO21D1 U3650 ( .A1(n965), .A2(n2148), .B(n2147), .Z(
        dp_cluster_1_mult_513_C418_n281) );
  XNR2D1 U3651 ( .A1(n1072), .A2(n1386), .ZN(n2047) );
  XNR2D1 U3652 ( .A1(n1072), .A2(n1385), .ZN(n2146) );
  XNR2D1 U3653 ( .A1(n1072), .A2(n1387), .ZN(n2048) );
  XNR2D1 U3654 ( .A1(n1072), .A2(n1390), .ZN(n2051) );
  XNR2D1 U3655 ( .A1(n1073), .A2(n1391), .ZN(n2052) );
  XNR2D1 U3656 ( .A1(n1072), .A2(n1392), .ZN(n2053) );
  XNR2D1 U3657 ( .A1(n1072), .A2(n1393), .ZN(n2054) );
  XNR2D1 U3658 ( .A1(n1072), .A2(n1394), .ZN(n2055) );
  XNR2D1 U3659 ( .A1(n1072), .A2(n1395), .ZN(n2056) );
  XNR2D1 U3660 ( .A1(n1072), .A2(n1396), .ZN(n2057) );
  XNR2D1 U3661 ( .A1(n1072), .A2(n1397), .ZN(n2058) );
  XNR2D1 U3662 ( .A1(n1072), .A2(n1398), .ZN(n2059) );
  XNR2D1 U3663 ( .A1(n1092), .A2(n1073), .ZN(n2060) );
  XNR2D1 U3664 ( .A1(s1_7_i[10]), .A2(W3_8_r[63]), .ZN(n2151) );
  AO21D1 U3665 ( .A1(n970), .A2(n2152), .B(n2151), .Z(
        dp_cluster_1_mult_513_C418_n296) );
  XNR2D1 U3666 ( .A1(n1075), .A2(n1386), .ZN(n2061) );
  XNR2D1 U3667 ( .A1(n1074), .A2(n1385), .ZN(n2150) );
  XNR2D1 U3668 ( .A1(n1074), .A2(n1387), .ZN(n2062) );
  XNR2D1 U3669 ( .A1(n1074), .A2(n1388), .ZN(n2063) );
  XNR2D1 U3670 ( .A1(n1074), .A2(n1389), .ZN(n2064) );
  XNR2D1 U3671 ( .A1(n1074), .A2(n1390), .ZN(n2065) );
  XNR2D1 U3672 ( .A1(n1075), .A2(n1391), .ZN(n2066) );
  XNR2D1 U3673 ( .A1(n1074), .A2(n1392), .ZN(n2067) );
  XNR2D1 U3674 ( .A1(n1074), .A2(n1393), .ZN(n2068) );
  XNR2D1 U3675 ( .A1(n1074), .A2(n1394), .ZN(n2069) );
  XNR2D1 U3676 ( .A1(n1074), .A2(n1395), .ZN(n2070) );
  XNR2D1 U3677 ( .A1(n1074), .A2(n1396), .ZN(n2071) );
  XNR2D1 U3678 ( .A1(n1074), .A2(n1397), .ZN(n2072) );
  XNR2D1 U3679 ( .A1(n1074), .A2(n1398), .ZN(n2073) );
  XNR2D1 U3680 ( .A1(n1092), .A2(n1076), .ZN(n2074) );
  XNR2D1 U3681 ( .A1(s1_7_i[8]), .A2(W3_8_r[63]), .ZN(n2075) );
  AO21D1 U3682 ( .A1(n968), .A2(n2092), .B(n2075), .Z(
        dp_cluster_1_mult_513_C418_n312) );
  XNR2D1 U3683 ( .A1(n1077), .A2(n1385), .ZN(n2076) );
  XNR2D1 U3684 ( .A1(n1077), .A2(n1386), .ZN(n2077) );
  XNR2D1 U3685 ( .A1(n1077), .A2(n1387), .ZN(n2078) );
  XNR2D1 U3686 ( .A1(n1077), .A2(n1388), .ZN(n2079) );
  XNR2D1 U3687 ( .A1(n1078), .A2(n1391), .ZN(n2082) );
  XNR2D1 U3688 ( .A1(n1077), .A2(n1392), .ZN(n2083) );
  XNR2D1 U3689 ( .A1(n1077), .A2(n1393), .ZN(n2084) );
  XNR2D1 U3690 ( .A1(n1077), .A2(n1394), .ZN(n2085) );
  XNR2D1 U3691 ( .A1(n1077), .A2(n1395), .ZN(n2086) );
  XNR2D1 U3692 ( .A1(n1077), .A2(n1396), .ZN(n2087) );
  XNR2D1 U3693 ( .A1(n1077), .A2(n1397), .ZN(n2088) );
  XNR2D1 U3694 ( .A1(n1077), .A2(n1398), .ZN(n2089) );
  XNR2D1 U3695 ( .A1(n1092), .A2(n1079), .ZN(n2091) );
  AO21D1 U3696 ( .A1(n966), .A2(n2110), .B(n2093), .Z(
        dp_cluster_1_mult_513_C418_n329) );
  XNR2D1 U3697 ( .A1(n1080), .A2(n1386), .ZN(n2095) );
  XNR2D1 U3698 ( .A1(n1080), .A2(n1387), .ZN(n2096) );
  XNR2D1 U3699 ( .A1(n1080), .A2(n1388), .ZN(n2097) );
  XNR2D1 U3700 ( .A1(n1080), .A2(n1389), .ZN(n2098) );
  XNR2D1 U3701 ( .A1(n1080), .A2(n1390), .ZN(n2099) );
  XNR2D1 U3702 ( .A1(n1081), .A2(n1391), .ZN(n2100) );
  XNR2D1 U3703 ( .A1(n1080), .A2(n1392), .ZN(n2101) );
  XNR2D1 U3704 ( .A1(n1080), .A2(n1393), .ZN(n2102) );
  XNR2D1 U3705 ( .A1(n1080), .A2(n1394), .ZN(n2103) );
  XNR2D1 U3706 ( .A1(n1080), .A2(n1395), .ZN(n2104) );
  XNR2D1 U3707 ( .A1(n1080), .A2(n1396), .ZN(n2105) );
  XNR2D1 U3708 ( .A1(n1080), .A2(n1397), .ZN(n2106) );
  XNR2D1 U3709 ( .A1(n1080), .A2(n1398), .ZN(n2107) );
  XNR2D1 U3710 ( .A1(n1092), .A2(n1082), .ZN(n2109) );
  AO21D1 U3711 ( .A1(n967), .A2(n2128), .B(n2111), .Z(
        dp_cluster_1_mult_513_C418_n345) );
  XNR2D1 U3712 ( .A1(n1083), .A2(n1386), .ZN(n2113) );
  XNR2D1 U3713 ( .A1(n1083), .A2(n1387), .ZN(n2114) );
  XNR2D1 U3714 ( .A1(n1083), .A2(n1388), .ZN(n2115) );
  XNR2D1 U3715 ( .A1(n1083), .A2(n1389), .ZN(n2116) );
  XNR2D1 U3716 ( .A1(n1083), .A2(n1390), .ZN(n2117) );
  XNR2D1 U3717 ( .A1(n1084), .A2(n1391), .ZN(n2118) );
  XNR2D1 U3718 ( .A1(n1083), .A2(n1392), .ZN(n2119) );
  XNR2D1 U3719 ( .A1(n1083), .A2(n1393), .ZN(n2120) );
  XNR2D1 U3720 ( .A1(n1083), .A2(n1394), .ZN(n2121) );
  XNR2D1 U3721 ( .A1(n1083), .A2(n1395), .ZN(n2122) );
  XNR2D1 U3722 ( .A1(n1083), .A2(n1396), .ZN(n2123) );
  XNR2D1 U3723 ( .A1(n1083), .A2(n1397), .ZN(n2124) );
  XNR2D1 U3724 ( .A1(n1083), .A2(n1398), .ZN(n2125) );
  XNR2D1 U3725 ( .A1(n1092), .A2(n1085), .ZN(n2127) );
  CKXOR2D1 U3726 ( .A1(n1102), .A2(W3_8_r[63]), .Z(n2129) );
  XNR2D1 U3727 ( .A1(n1102), .A2(W3_8_r[62]), .ZN(n2130) );
  MOAI22D1 U3728 ( .A1(n2130), .A2(n2144), .B1(n2129), .B2(s1_7_i[1]), .ZN(
        dp_cluster_1_mult_513_C418_n362) );
  XNR2D1 U3729 ( .A1(n1101), .A2(W3_8_r[61]), .ZN(n2131) );
  XNR2D1 U3730 ( .A1(n1101), .A2(W3_8_r[60]), .ZN(n2132) );
  XNR2D1 U3731 ( .A1(n1101), .A2(W3_8_r[59]), .ZN(n2133) );
  XNR2D1 U3732 ( .A1(n1101), .A2(W3_8_r[58]), .ZN(n2134) );
  XNR2D1 U3733 ( .A1(n1101), .A2(W3_8_r[57]), .ZN(n2135) );
  XNR2D1 U3734 ( .A1(n1101), .A2(W3_8_r[56]), .ZN(n2136) );
  XNR2D1 U3735 ( .A1(n1101), .A2(W3_8_r[55]), .ZN(n2137) );
  XNR2D1 U3736 ( .A1(n1101), .A2(W3_8_r[54]), .ZN(n2138) );
  XNR2D1 U3737 ( .A1(n1101), .A2(W3_8_r[53]), .ZN(n2139) );
  XNR2D1 U3738 ( .A1(n1101), .A2(W3_8_r[52]), .ZN(n2140) );
  XNR2D1 U3739 ( .A1(n1101), .A2(W3_8_r[51]), .ZN(n2141) );
  XNR2D1 U3740 ( .A1(n1101), .A2(W3_8_r[50]), .ZN(n2142) );
  XNR2D1 U3741 ( .A1(n1102), .A2(W3_8_r[49]), .ZN(n2143) );
  XNR2D1 U3742 ( .A1(W3_8_r[61]), .A2(s1_7_i[16]), .ZN(n2156) );
  XNR2D1 U3743 ( .A1(s1_7_i[14]), .A2(W3_8_r[63]), .ZN(n2157) );
  XNR2D1 U3744 ( .A1(n1029), .A2(n1419), .ZN(n2202) );
  XNR2D1 U3745 ( .A1(n1029), .A2(s1_7_r[11]), .ZN(n2164) );
  XNR2D1 U3746 ( .A1(n1028), .A2(n1418), .ZN(n2201) );
  XNR2D1 U3747 ( .A1(s1_7_r[6]), .A2(W3_8_i[63]), .ZN(n2245) );
  XNR2D1 U3748 ( .A1(n1037), .A2(n1415), .ZN(n2246) );
  XNR2D1 U3749 ( .A1(n1037), .A2(s1_7_r[5]), .ZN(n2165) );
  XNR2D1 U3750 ( .A1(s1_7_r[4]), .A2(W3_8_i[63]), .ZN(n2263) );
  XNR2D1 U3751 ( .A1(n1040), .A2(n1415), .ZN(n2264) );
  XNR2D1 U3752 ( .A1(n1040), .A2(s1_7_r[3]), .ZN(n2166) );
  XNR2D1 U3753 ( .A1(n1034), .A2(n1420), .ZN(n2233) );
  XNR2D1 U3754 ( .A1(n1034), .A2(s1_7_r[7]), .ZN(n2167) );
  XNR2D1 U3755 ( .A1(n1034), .A2(n1419), .ZN(n2232) );
  XNR2D1 U3756 ( .A1(n1026), .A2(n1426), .ZN(n2195) );
  XNR2D1 U3757 ( .A1(n1026), .A2(s1_7_r[13]), .ZN(n2168) );
  XNR2D1 U3758 ( .A1(n1026), .A2(n1425), .ZN(n2194) );
  XNR2D1 U3759 ( .A1(n2170), .A2(n2169), .ZN(dp_cluster_1_mult_512_C418_n162)
         );
  XNR2D1 U3760 ( .A1(n1023), .A2(s1_7_r[15]), .ZN(n2171) );
  XNR2D1 U3761 ( .A1(n1031), .A2(s1_7_r[9]), .ZN(n2172) );
  XNR2D1 U3762 ( .A1(n1023), .A2(n1418), .ZN(n2173) );
  XNR2D1 U3763 ( .A1(s1_7_r[16]), .A2(W3_8_i[60]), .ZN(n2305) );
  XNR2D1 U3764 ( .A1(n1023), .A2(n1419), .ZN(n2174) );
  XNR2D1 U3765 ( .A1(n1023), .A2(n1420), .ZN(n2175) );
  XNR2D1 U3766 ( .A1(n1023), .A2(n1421), .ZN(n2176) );
  XNR2D1 U3767 ( .A1(n1023), .A2(n1422), .ZN(n2177) );
  XNR2D1 U3768 ( .A1(n1023), .A2(n1423), .ZN(n2178) );
  XNR2D1 U3769 ( .A1(n1023), .A2(n1424), .ZN(n2179) );
  XNR2D1 U3770 ( .A1(n1023), .A2(n1425), .ZN(n2180) );
  XNR2D1 U3771 ( .A1(n1023), .A2(n1426), .ZN(n2181) );
  XNR2D1 U3772 ( .A1(n1023), .A2(n1427), .ZN(n2182) );
  XNR2D1 U3773 ( .A1(n1023), .A2(n1428), .ZN(n2183) );
  XNR2D1 U3774 ( .A1(n1099), .A2(n1024), .ZN(n2184) );
  XNR2D1 U3775 ( .A1(n1025), .A2(n1416), .ZN(n2185) );
  XNR2D1 U3776 ( .A1(n1025), .A2(n1415), .ZN(n2312) );
  XNR2D1 U3777 ( .A1(n1025), .A2(n1417), .ZN(n2186) );
  XNR2D1 U3778 ( .A1(n1025), .A2(n1418), .ZN(n2187) );
  XNR2D1 U3779 ( .A1(n1026), .A2(n1419), .ZN(n2188) );
  XNR2D1 U3780 ( .A1(n1025), .A2(n1420), .ZN(n2189) );
  XNR2D1 U3781 ( .A1(n1025), .A2(n1421), .ZN(n2190) );
  XNR2D1 U3782 ( .A1(n1025), .A2(n1422), .ZN(n2191) );
  XNR2D1 U3783 ( .A1(n1025), .A2(n1423), .ZN(n2192) );
  XNR2D1 U3784 ( .A1(n1025), .A2(n1424), .ZN(n2193) );
  XNR2D1 U3785 ( .A1(n1025), .A2(n1427), .ZN(n2196) );
  XNR2D1 U3786 ( .A1(n1025), .A2(n1428), .ZN(n2197) );
  XNR2D1 U3787 ( .A1(n1098), .A2(n1027), .ZN(n2198) );
  XNR2D1 U3788 ( .A1(s1_7_r[12]), .A2(W3_8_i[63]), .ZN(n2299) );
  AO21D1 U3789 ( .A1(n971), .A2(n2300), .B(n2299), .Z(
        dp_cluster_1_mult_512_C418_n281) );
  XNR2D1 U3790 ( .A1(n1028), .A2(n1416), .ZN(n2199) );
  XNR2D1 U3791 ( .A1(n1028), .A2(n1415), .ZN(n2298) );
  XNR2D1 U3792 ( .A1(n1028), .A2(n1417), .ZN(n2200) );
  XNR2D1 U3793 ( .A1(n1028), .A2(n1420), .ZN(n2203) );
  XNR2D1 U3794 ( .A1(n1029), .A2(n1421), .ZN(n2204) );
  XNR2D1 U3795 ( .A1(n1028), .A2(n1422), .ZN(n2205) );
  XNR2D1 U3796 ( .A1(n1028), .A2(n1423), .ZN(n2206) );
  XNR2D1 U3797 ( .A1(n1028), .A2(n1424), .ZN(n2207) );
  XNR2D1 U3798 ( .A1(n1028), .A2(n1425), .ZN(n2208) );
  XNR2D1 U3799 ( .A1(n1028), .A2(n1426), .ZN(n2209) );
  XNR2D1 U3800 ( .A1(n1028), .A2(n1427), .ZN(n2210) );
  XNR2D1 U3801 ( .A1(n1028), .A2(n1428), .ZN(n2211) );
  XNR2D1 U3802 ( .A1(n1098), .A2(n1029), .ZN(n2212) );
  XNR2D1 U3803 ( .A1(s1_7_r[10]), .A2(W3_8_i[63]), .ZN(n2303) );
  AO21D1 U3804 ( .A1(n976), .A2(n2304), .B(n2303), .Z(
        dp_cluster_1_mult_512_C418_n296) );
  XNR2D1 U3805 ( .A1(n1031), .A2(n1416), .ZN(n2213) );
  XNR2D1 U3806 ( .A1(n1030), .A2(n1415), .ZN(n2302) );
  XNR2D1 U3807 ( .A1(n1030), .A2(n1417), .ZN(n2214) );
  XNR2D1 U3808 ( .A1(n1030), .A2(n1418), .ZN(n2215) );
  XNR2D1 U3809 ( .A1(n1030), .A2(n1419), .ZN(n2216) );
  XNR2D1 U3810 ( .A1(n1030), .A2(n1420), .ZN(n2217) );
  XNR2D1 U3811 ( .A1(n1031), .A2(n1421), .ZN(n2218) );
  XNR2D1 U3812 ( .A1(n1030), .A2(n1422), .ZN(n2219) );
  XNR2D1 U3813 ( .A1(n1030), .A2(n1423), .ZN(n2220) );
  XNR2D1 U3814 ( .A1(n1030), .A2(n1424), .ZN(n2221) );
  XNR2D1 U3815 ( .A1(n1030), .A2(n1425), .ZN(n2222) );
  XNR2D1 U3816 ( .A1(n1030), .A2(n1426), .ZN(n2223) );
  XNR2D1 U3817 ( .A1(n1030), .A2(n1427), .ZN(n2224) );
  XNR2D1 U3818 ( .A1(n1030), .A2(n1428), .ZN(n2225) );
  XNR2D1 U3819 ( .A1(n1098), .A2(n1032), .ZN(n2226) );
  XNR2D1 U3820 ( .A1(s1_7_r[8]), .A2(W3_8_i[63]), .ZN(n2227) );
  AO21D1 U3821 ( .A1(n974), .A2(n2244), .B(n2227), .Z(
        dp_cluster_1_mult_512_C418_n312) );
  XNR2D1 U3822 ( .A1(n1033), .A2(n1415), .ZN(n2228) );
  XNR2D1 U3823 ( .A1(n1033), .A2(n1416), .ZN(n2229) );
  XNR2D1 U3824 ( .A1(n1033), .A2(n1417), .ZN(n2230) );
  XNR2D1 U3825 ( .A1(n1033), .A2(n1418), .ZN(n2231) );
  XNR2D1 U3826 ( .A1(n1034), .A2(n1421), .ZN(n2234) );
  XNR2D1 U3827 ( .A1(n1033), .A2(n1422), .ZN(n2235) );
  XNR2D1 U3828 ( .A1(n1033), .A2(n1423), .ZN(n2236) );
  XNR2D1 U3829 ( .A1(n1033), .A2(n1424), .ZN(n2237) );
  XNR2D1 U3830 ( .A1(n1033), .A2(n1425), .ZN(n2238) );
  XNR2D1 U3831 ( .A1(n1033), .A2(n1426), .ZN(n2239) );
  XNR2D1 U3832 ( .A1(n1033), .A2(n1427), .ZN(n2240) );
  XNR2D1 U3833 ( .A1(n1033), .A2(n1428), .ZN(n2241) );
  XNR2D1 U3834 ( .A1(n1098), .A2(n1035), .ZN(n2243) );
  AO21D1 U3835 ( .A1(n972), .A2(n2262), .B(n2245), .Z(
        dp_cluster_1_mult_512_C418_n329) );
  XNR2D1 U3836 ( .A1(n1036), .A2(n1416), .ZN(n2247) );
  XNR2D1 U3837 ( .A1(n1036), .A2(n1417), .ZN(n2248) );
  XNR2D1 U3838 ( .A1(n1036), .A2(n1418), .ZN(n2249) );
  XNR2D1 U3839 ( .A1(n1036), .A2(n1419), .ZN(n2250) );
  XNR2D1 U3840 ( .A1(n1036), .A2(n1420), .ZN(n2251) );
  XNR2D1 U3841 ( .A1(n1037), .A2(n1421), .ZN(n2252) );
  XNR2D1 U3842 ( .A1(n1036), .A2(n1422), .ZN(n2253) );
  XNR2D1 U3843 ( .A1(n1036), .A2(n1423), .ZN(n2254) );
  XNR2D1 U3844 ( .A1(n1036), .A2(n1424), .ZN(n2255) );
  XNR2D1 U3845 ( .A1(n1036), .A2(n1425), .ZN(n2256) );
  XNR2D1 U3846 ( .A1(n1036), .A2(n1426), .ZN(n2257) );
  XNR2D1 U3847 ( .A1(n1036), .A2(n1427), .ZN(n2258) );
  XNR2D1 U3848 ( .A1(n1036), .A2(n1428), .ZN(n2259) );
  XNR2D1 U3849 ( .A1(n1098), .A2(n1038), .ZN(n2261) );
  AO21D1 U3850 ( .A1(n973), .A2(n2280), .B(n2263), .Z(
        dp_cluster_1_mult_512_C418_n345) );
  XNR2D1 U3851 ( .A1(n1039), .A2(n1416), .ZN(n2265) );
  XNR2D1 U3852 ( .A1(n1039), .A2(n1417), .ZN(n2266) );
  XNR2D1 U3853 ( .A1(n1039), .A2(n1418), .ZN(n2267) );
  XNR2D1 U3854 ( .A1(n1039), .A2(n1419), .ZN(n2268) );
  XNR2D1 U3855 ( .A1(n1039), .A2(n1420), .ZN(n2269) );
  XNR2D1 U3856 ( .A1(n1040), .A2(n1421), .ZN(n2270) );
  XNR2D1 U3857 ( .A1(n1039), .A2(n1422), .ZN(n2271) );
  XNR2D1 U3858 ( .A1(n1039), .A2(n1423), .ZN(n2272) );
  XNR2D1 U3859 ( .A1(n1039), .A2(n1424), .ZN(n2273) );
  XNR2D1 U3860 ( .A1(n1039), .A2(n1425), .ZN(n2274) );
  XNR2D1 U3861 ( .A1(n1039), .A2(n1426), .ZN(n2275) );
  XNR2D1 U3862 ( .A1(n1039), .A2(n1427), .ZN(n2276) );
  XNR2D1 U3863 ( .A1(n1039), .A2(n1428), .ZN(n2277) );
  XNR2D1 U3864 ( .A1(n1098), .A2(n1041), .ZN(n2279) );
  CKXOR2D1 U3865 ( .A1(n1108), .A2(W3_8_i[63]), .Z(n2281) );
  XNR2D1 U3866 ( .A1(n1108), .A2(W3_8_i[62]), .ZN(n2282) );
  MOAI22D1 U3867 ( .A1(n2282), .A2(n2296), .B1(n2281), .B2(s1_7_r[1]), .ZN(
        dp_cluster_1_mult_512_C418_n362) );
  XNR2D1 U3868 ( .A1(n1107), .A2(W3_8_i[61]), .ZN(n2283) );
  XNR2D1 U3869 ( .A1(n1107), .A2(W3_8_i[60]), .ZN(n2284) );
  XNR2D1 U3870 ( .A1(n1107), .A2(W3_8_i[59]), .ZN(n2285) );
  XNR2D1 U3871 ( .A1(n1107), .A2(W3_8_i[58]), .ZN(n2286) );
  XNR2D1 U3872 ( .A1(n1107), .A2(W3_8_i[57]), .ZN(n2287) );
  XNR2D1 U3873 ( .A1(n1107), .A2(W3_8_i[56]), .ZN(n2288) );
  XNR2D1 U3874 ( .A1(n1107), .A2(W3_8_i[55]), .ZN(n2289) );
  XNR2D1 U3875 ( .A1(n1107), .A2(W3_8_i[54]), .ZN(n2290) );
  XNR2D1 U3876 ( .A1(n1107), .A2(W3_8_i[53]), .ZN(n2291) );
  XNR2D1 U3877 ( .A1(n1107), .A2(W3_8_i[52]), .ZN(n2292) );
  XNR2D1 U3878 ( .A1(n1107), .A2(W3_8_i[51]), .ZN(n2293) );
  XNR2D1 U3879 ( .A1(n1107), .A2(W3_8_i[50]), .ZN(n2294) );
  XNR2D1 U3880 ( .A1(n1108), .A2(W3_8_i[49]), .ZN(n2295) );
  XNR2D1 U3881 ( .A1(W3_8_i[61]), .A2(s1_7_r[16]), .ZN(n2308) );
  XNR2D1 U3882 ( .A1(s1_7_r[14]), .A2(W3_8_i[63]), .ZN(n2309) );
  XNR2D1 U3883 ( .A1(n1050), .A2(n1404), .ZN(n2375) );
  XNR2D1 U3884 ( .A1(n1051), .A2(s1_5_i[11]), .ZN(n2337) );
  XNR2D1 U3885 ( .A1(n1051), .A2(n1403), .ZN(n2374) );
  XNR2D1 U3886 ( .A1(s1_5_i[6]), .A2(W1_8_i[63]), .ZN(n2418) );
  XNR2D1 U3887 ( .A1(n1058), .A2(n1400), .ZN(n2419) );
  XNR2D1 U3888 ( .A1(n1059), .A2(s1_5_i[5]), .ZN(n2338) );
  XNR2D1 U3889 ( .A1(s1_5_i[4]), .A2(W1_8_i[63]), .ZN(n2436) );
  XNR2D1 U3890 ( .A1(n1062), .A2(n1400), .ZN(n2437) );
  XNR2D1 U3891 ( .A1(n1063), .A2(s1_5_i[3]), .ZN(n2339) );
  XNR2D1 U3892 ( .A1(n1055), .A2(n1405), .ZN(n2406) );
  XNR2D1 U3893 ( .A1(n1056), .A2(s1_5_i[7]), .ZN(n2340) );
  XNR2D1 U3894 ( .A1(n1057), .A2(n1404), .ZN(n2405) );
  XNR2D1 U3895 ( .A1(n1047), .A2(n1411), .ZN(n2368) );
  XNR2D1 U3896 ( .A1(n1048), .A2(s1_5_i[13]), .ZN(n2341) );
  XNR2D1 U3897 ( .A1(n1049), .A2(n1410), .ZN(n2367) );
  XNR2D1 U3898 ( .A1(n2343), .A2(n2342), .ZN(dp_cluster_2_mult_486_C409_n162)
         );
  XNR2D1 U3899 ( .A1(n1045), .A2(s1_5_i[15]), .ZN(n2344) );
  XNR2D1 U3900 ( .A1(n1053), .A2(s1_5_i[9]), .ZN(n2345) );
  XNR2D1 U3901 ( .A1(n1046), .A2(n1403), .ZN(n2346) );
  XNR2D1 U3902 ( .A1(s1_5_i[16]), .A2(W1_8_i[60]), .ZN(n2478) );
  XNR2D1 U3903 ( .A1(n1046), .A2(n1404), .ZN(n2347) );
  XNR2D1 U3904 ( .A1(n1046), .A2(n1405), .ZN(n2348) );
  XNR2D1 U3905 ( .A1(n1046), .A2(n1406), .ZN(n2349) );
  XNR2D1 U3906 ( .A1(n1046), .A2(n1407), .ZN(n2350) );
  XNR2D1 U3907 ( .A1(n1046), .A2(n1408), .ZN(n2351) );
  XNR2D1 U3908 ( .A1(n1046), .A2(n1409), .ZN(n2352) );
  XNR2D1 U3909 ( .A1(n1046), .A2(n1410), .ZN(n2353) );
  XNR2D1 U3910 ( .A1(n1046), .A2(n1411), .ZN(n2354) );
  XNR2D1 U3911 ( .A1(n1046), .A2(n1412), .ZN(n2355) );
  XNR2D1 U3912 ( .A1(n1046), .A2(n1413), .ZN(n2356) );
  XNR2D1 U3913 ( .A1(n1097), .A2(n1046), .ZN(n2357) );
  XNR2D1 U3914 ( .A1(n1048), .A2(n1401), .ZN(n2358) );
  XNR2D1 U3915 ( .A1(n1048), .A2(n1400), .ZN(n2485) );
  XNR2D1 U3916 ( .A1(n1048), .A2(n1402), .ZN(n2359) );
  XNR2D1 U3917 ( .A1(n1048), .A2(n1403), .ZN(n2360) );
  XNR2D1 U3918 ( .A1(n1048), .A2(n1404), .ZN(n2361) );
  XNR2D1 U3919 ( .A1(n1048), .A2(n1405), .ZN(n2362) );
  XNR2D1 U3920 ( .A1(n1048), .A2(n1406), .ZN(n2363) );
  XNR2D1 U3921 ( .A1(n1048), .A2(n1407), .ZN(n2364) );
  XNR2D1 U3922 ( .A1(n1048), .A2(n1408), .ZN(n2365) );
  XNR2D1 U3923 ( .A1(n1048), .A2(n1409), .ZN(n2366) );
  XNR2D1 U3924 ( .A1(n1048), .A2(n1412), .ZN(n2369) );
  XNR2D1 U3925 ( .A1(n1048), .A2(n1413), .ZN(n2370) );
  XNR2D1 U3926 ( .A1(n1097), .A2(n1049), .ZN(n2371) );
  XNR2D1 U3927 ( .A1(s1_5_i[12]), .A2(W1_8_i[63]), .ZN(n2472) );
  AO21D1 U3928 ( .A1(n977), .A2(n2473), .B(n2472), .Z(
        dp_cluster_2_mult_486_C409_n281) );
  XNR2D1 U3929 ( .A1(n1051), .A2(n1401), .ZN(n2372) );
  XNR2D1 U3930 ( .A1(n1051), .A2(n1400), .ZN(n2471) );
  XNR2D1 U3931 ( .A1(n1051), .A2(n1402), .ZN(n2373) );
  XNR2D1 U3932 ( .A1(n1051), .A2(n1405), .ZN(n2376) );
  XNR2D1 U3933 ( .A1(n1051), .A2(n1406), .ZN(n2377) );
  XNR2D1 U3934 ( .A1(n1051), .A2(n1407), .ZN(n2378) );
  XNR2D1 U3935 ( .A1(n1051), .A2(n1408), .ZN(n2379) );
  XNR2D1 U3936 ( .A1(n1051), .A2(n1409), .ZN(n2380) );
  XNR2D1 U3937 ( .A1(n1051), .A2(n1410), .ZN(n2381) );
  XNR2D1 U3938 ( .A1(n1051), .A2(n1411), .ZN(n2382) );
  XNR2D1 U3939 ( .A1(n1051), .A2(n1412), .ZN(n2383) );
  XNR2D1 U3940 ( .A1(n1051), .A2(n1413), .ZN(n2384) );
  XNR2D1 U3941 ( .A1(n1097), .A2(n1051), .ZN(n2385) );
  XNR2D1 U3942 ( .A1(s1_5_i[10]), .A2(W1_8_i[63]), .ZN(n2476) );
  AO21D1 U3943 ( .A1(n982), .A2(n2477), .B(n2476), .Z(
        dp_cluster_2_mult_486_C409_n296) );
  XNR2D1 U3944 ( .A1(n1054), .A2(n1401), .ZN(n2386) );
  XNR2D1 U3945 ( .A1(n1053), .A2(n1400), .ZN(n2475) );
  XNR2D1 U3946 ( .A1(n1053), .A2(n1402), .ZN(n2387) );
  XNR2D1 U3947 ( .A1(n1053), .A2(n1403), .ZN(n2388) );
  XNR2D1 U3948 ( .A1(n1053), .A2(n1404), .ZN(n2389) );
  XNR2D1 U3949 ( .A1(n1053), .A2(n1405), .ZN(n2390) );
  XNR2D1 U3950 ( .A1(n1053), .A2(n1406), .ZN(n2391) );
  XNR2D1 U3951 ( .A1(n1053), .A2(n1407), .ZN(n2392) );
  XNR2D1 U3952 ( .A1(n1053), .A2(n1408), .ZN(n2393) );
  XNR2D1 U3953 ( .A1(n1053), .A2(n1409), .ZN(n2394) );
  XNR2D1 U3954 ( .A1(n1053), .A2(n1410), .ZN(n2395) );
  XNR2D1 U3955 ( .A1(n1053), .A2(n1411), .ZN(n2396) );
  XNR2D1 U3956 ( .A1(n1053), .A2(n1412), .ZN(n2397) );
  XNR2D1 U3957 ( .A1(n1053), .A2(n1413), .ZN(n2398) );
  XNR2D1 U3958 ( .A1(n1097), .A2(n1054), .ZN(n2399) );
  XNR2D1 U3959 ( .A1(s1_5_i[8]), .A2(W1_8_i[63]), .ZN(n2400) );
  AO21D1 U3960 ( .A1(n980), .A2(n2417), .B(n2400), .Z(
        dp_cluster_2_mult_486_C409_n312) );
  XNR2D1 U3961 ( .A1(n1056), .A2(n1400), .ZN(n2401) );
  XNR2D1 U3962 ( .A1(n1056), .A2(n1401), .ZN(n2402) );
  XNR2D1 U3963 ( .A1(n1056), .A2(n1402), .ZN(n2403) );
  XNR2D1 U3964 ( .A1(n1056), .A2(n1403), .ZN(n2404) );
  XNR2D1 U3965 ( .A1(n1056), .A2(n1406), .ZN(n2407) );
  XNR2D1 U3966 ( .A1(n1056), .A2(n1407), .ZN(n2408) );
  XNR2D1 U3967 ( .A1(n1056), .A2(n1408), .ZN(n2409) );
  XNR2D1 U3968 ( .A1(n1056), .A2(n1409), .ZN(n2410) );
  XNR2D1 U3969 ( .A1(n1056), .A2(n1410), .ZN(n2411) );
  XNR2D1 U3970 ( .A1(n1056), .A2(n1411), .ZN(n2412) );
  XNR2D1 U3971 ( .A1(n1056), .A2(n1412), .ZN(n2413) );
  XNR2D1 U3972 ( .A1(n1056), .A2(n1413), .ZN(n2414) );
  XNR2D1 U3973 ( .A1(n1096), .A2(n1057), .ZN(n2416) );
  AO21D1 U3974 ( .A1(n978), .A2(n2435), .B(n2418), .Z(
        dp_cluster_2_mult_486_C409_n329) );
  XNR2D1 U3975 ( .A1(n1059), .A2(n1401), .ZN(n2420) );
  XNR2D1 U3976 ( .A1(n1059), .A2(n1402), .ZN(n2421) );
  XNR2D1 U3977 ( .A1(n1059), .A2(n1403), .ZN(n2422) );
  XNR2D1 U3978 ( .A1(n1059), .A2(n1404), .ZN(n2423) );
  XNR2D1 U3979 ( .A1(n1059), .A2(n1405), .ZN(n2424) );
  XNR2D1 U3980 ( .A1(n1059), .A2(n1406), .ZN(n2425) );
  XNR2D1 U3981 ( .A1(n1059), .A2(n1407), .ZN(n2426) );
  XNR2D1 U3982 ( .A1(n1059), .A2(n1408), .ZN(n2427) );
  XNR2D1 U3983 ( .A1(n1059), .A2(n1409), .ZN(n2428) );
  XNR2D1 U3984 ( .A1(n1059), .A2(n1410), .ZN(n2429) );
  XNR2D1 U3985 ( .A1(n1059), .A2(n1411), .ZN(n2430) );
  XNR2D1 U3986 ( .A1(n1059), .A2(n1412), .ZN(n2431) );
  XNR2D1 U3987 ( .A1(n1059), .A2(n1413), .ZN(n2432) );
  XNR2D1 U3988 ( .A1(n1096), .A2(n1060), .ZN(n2434) );
  AO21D1 U3989 ( .A1(n979), .A2(n2453), .B(n2436), .Z(
        dp_cluster_2_mult_486_C409_n345) );
  XNR2D1 U3990 ( .A1(n1062), .A2(n1401), .ZN(n2438) );
  XNR2D1 U3991 ( .A1(n1062), .A2(n1402), .ZN(n2439) );
  XNR2D1 U3992 ( .A1(n1062), .A2(n1403), .ZN(n2440) );
  XNR2D1 U3993 ( .A1(n1062), .A2(n1404), .ZN(n2441) );
  XNR2D1 U3994 ( .A1(n1062), .A2(n1405), .ZN(n2442) );
  XNR2D1 U3995 ( .A1(n1062), .A2(n1406), .ZN(n2443) );
  XNR2D1 U3996 ( .A1(n1062), .A2(n1407), .ZN(n2444) );
  XNR2D1 U3997 ( .A1(n1062), .A2(n1408), .ZN(n2445) );
  XNR2D1 U3998 ( .A1(n1062), .A2(n1409), .ZN(n2446) );
  XNR2D1 U3999 ( .A1(n1062), .A2(n1410), .ZN(n2447) );
  XNR2D1 U4000 ( .A1(n1062), .A2(n1411), .ZN(n2448) );
  XNR2D1 U4001 ( .A1(n1062), .A2(n1412), .ZN(n2449) );
  XNR2D1 U4002 ( .A1(n1062), .A2(n1413), .ZN(n2450) );
  XNR2D1 U4003 ( .A1(n1096), .A2(n1063), .ZN(n2452) );
  CKXOR2D1 U4004 ( .A1(n1106), .A2(W1_8_i[63]), .Z(n2454) );
  XNR2D1 U4005 ( .A1(n1106), .A2(W1_8_i[62]), .ZN(n2455) );
  MOAI22D1 U4006 ( .A1(n2455), .A2(n2469), .B1(n2454), .B2(s1_5_i[1]), .ZN(
        dp_cluster_2_mult_486_C409_n362) );
  XNR2D1 U4007 ( .A1(n1105), .A2(W1_8_i[61]), .ZN(n2456) );
  XNR2D1 U4008 ( .A1(n1106), .A2(W1_8_i[60]), .ZN(n2457) );
  XNR2D1 U4009 ( .A1(n1106), .A2(W1_8_i[59]), .ZN(n2458) );
  XNR2D1 U4010 ( .A1(n1105), .A2(W1_8_i[58]), .ZN(n2459) );
  XNR2D1 U4011 ( .A1(n1105), .A2(W1_8_i[57]), .ZN(n2460) );
  XNR2D1 U4012 ( .A1(n1105), .A2(W1_8_i[56]), .ZN(n2461) );
  XNR2D1 U4013 ( .A1(n1105), .A2(W1_8_i[55]), .ZN(n2462) );
  XNR2D1 U4014 ( .A1(n1105), .A2(W1_8_i[54]), .ZN(n2463) );
  XNR2D1 U4015 ( .A1(n1105), .A2(W1_8_i[53]), .ZN(n2464) );
  XNR2D1 U4016 ( .A1(n1105), .A2(W1_8_i[52]), .ZN(n2465) );
  XNR2D1 U4017 ( .A1(n1105), .A2(W1_8_i[51]), .ZN(n2466) );
  XNR2D1 U4018 ( .A1(n1105), .A2(W1_8_i[50]), .ZN(n2467) );
  XNR2D1 U4019 ( .A1(n1105), .A2(W1_8_i[49]), .ZN(n2468) );
  XNR2D1 U4020 ( .A1(W1_8_i[61]), .A2(s1_5_i[16]), .ZN(n2481) );
  XNR2D1 U4021 ( .A1(s1_5_i[14]), .A2(W1_8_i[63]), .ZN(n2482) );
  XNR2D1 U4022 ( .A1(n1006), .A2(n1374), .ZN(n2527) );
  XNR2D1 U4023 ( .A1(n1007), .A2(s1_5_r[11]), .ZN(n2489) );
  XNR2D1 U4024 ( .A1(n1007), .A2(n1373), .ZN(n2526) );
  XNR2D1 U4025 ( .A1(s1_5_r[6]), .A2(W1_8_r[63]), .ZN(n2570) );
  XNR2D1 U4026 ( .A1(n1014), .A2(n1370), .ZN(n2571) );
  XNR2D1 U4027 ( .A1(n1015), .A2(s1_5_r[5]), .ZN(n2490) );
  XNR2D1 U4028 ( .A1(s1_5_r[4]), .A2(W1_8_r[63]), .ZN(n2588) );
  XNR2D1 U4029 ( .A1(n1018), .A2(n1370), .ZN(n2589) );
  XNR2D1 U4030 ( .A1(n1019), .A2(s1_5_r[3]), .ZN(n2491) );
  XNR2D1 U4031 ( .A1(n1011), .A2(n1375), .ZN(n2558) );
  XNR2D1 U4032 ( .A1(n1012), .A2(s1_5_r[7]), .ZN(n2492) );
  XNR2D1 U4033 ( .A1(n1013), .A2(n1374), .ZN(n2557) );
  XNR2D1 U4034 ( .A1(n1003), .A2(n1381), .ZN(n2520) );
  XNR2D1 U4035 ( .A1(n1004), .A2(s1_5_r[13]), .ZN(n2493) );
  XNR2D1 U4036 ( .A1(n1005), .A2(n1380), .ZN(n2519) );
  XNR2D1 U4037 ( .A1(n2495), .A2(n2494), .ZN(dp_cluster_2_mult_485_C409_n162)
         );
  XNR2D1 U4038 ( .A1(n1001), .A2(s1_5_r[15]), .ZN(n2496) );
  XNR2D1 U4039 ( .A1(n1009), .A2(s1_5_r[9]), .ZN(n2497) );
  XNR2D1 U4040 ( .A1(n1002), .A2(n1373), .ZN(n2498) );
  XNR2D1 U4041 ( .A1(s1_5_r[16]), .A2(W1_8_r[60]), .ZN(n2630) );
  XNR2D1 U4042 ( .A1(n1002), .A2(n1374), .ZN(n2499) );
  XNR2D1 U4043 ( .A1(n1002), .A2(n1375), .ZN(n2500) );
  XNR2D1 U4044 ( .A1(n1002), .A2(n1376), .ZN(n2501) );
  XNR2D1 U4045 ( .A1(n1002), .A2(n1377), .ZN(n2502) );
  XNR2D1 U4046 ( .A1(n1002), .A2(n1378), .ZN(n2503) );
  XNR2D1 U4047 ( .A1(n1002), .A2(n1379), .ZN(n2504) );
  XNR2D1 U4048 ( .A1(n1002), .A2(n1380), .ZN(n2505) );
  XNR2D1 U4049 ( .A1(n1002), .A2(n1381), .ZN(n2506) );
  XNR2D1 U4050 ( .A1(n1002), .A2(n1382), .ZN(n2507) );
  XNR2D1 U4051 ( .A1(n1002), .A2(n1383), .ZN(n2508) );
  XNR2D1 U4052 ( .A1(n1091), .A2(n1002), .ZN(n2509) );
  XNR2D1 U4053 ( .A1(n1004), .A2(n1371), .ZN(n2510) );
  XNR2D1 U4054 ( .A1(n1004), .A2(n1370), .ZN(n2637) );
  XNR2D1 U4055 ( .A1(n1004), .A2(n1372), .ZN(n2511) );
  XNR2D1 U4056 ( .A1(n1004), .A2(n1373), .ZN(n2512) );
  XNR2D1 U4057 ( .A1(n1004), .A2(n1374), .ZN(n2513) );
  XNR2D1 U4058 ( .A1(n1004), .A2(n1375), .ZN(n2514) );
  XNR2D1 U4059 ( .A1(n1004), .A2(n1376), .ZN(n2515) );
  XNR2D1 U4060 ( .A1(n1004), .A2(n1377), .ZN(n2516) );
  XNR2D1 U4061 ( .A1(n1004), .A2(n1378), .ZN(n2517) );
  XNR2D1 U4062 ( .A1(n1004), .A2(n1379), .ZN(n2518) );
  XNR2D1 U4063 ( .A1(n1004), .A2(n1382), .ZN(n2521) );
  XNR2D1 U4064 ( .A1(n1004), .A2(n1383), .ZN(n2522) );
  XNR2D1 U4065 ( .A1(n1091), .A2(n1005), .ZN(n2523) );
  XNR2D1 U4066 ( .A1(s1_5_r[12]), .A2(W1_8_r[63]), .ZN(n2624) );
  AO21D1 U4067 ( .A1(n983), .A2(n2625), .B(n2624), .Z(
        dp_cluster_2_mult_485_C409_n281) );
  XNR2D1 U4068 ( .A1(n1007), .A2(n1371), .ZN(n2524) );
  XNR2D1 U4069 ( .A1(n1007), .A2(n1370), .ZN(n2623) );
  XNR2D1 U4070 ( .A1(n1007), .A2(n1372), .ZN(n2525) );
  XNR2D1 U4071 ( .A1(n1007), .A2(n1375), .ZN(n2528) );
  XNR2D1 U4072 ( .A1(n1007), .A2(n1376), .ZN(n2529) );
  XNR2D1 U4073 ( .A1(n1007), .A2(n1377), .ZN(n2530) );
  XNR2D1 U4074 ( .A1(n1007), .A2(n1378), .ZN(n2531) );
  XNR2D1 U4075 ( .A1(n1007), .A2(n1379), .ZN(n2532) );
  XNR2D1 U4076 ( .A1(n1007), .A2(n1380), .ZN(n2533) );
  XNR2D1 U4077 ( .A1(n1007), .A2(n1381), .ZN(n2534) );
  XNR2D1 U4078 ( .A1(n1007), .A2(n1382), .ZN(n2535) );
  XNR2D1 U4079 ( .A1(n1007), .A2(n1383), .ZN(n2536) );
  XNR2D1 U4080 ( .A1(n1091), .A2(n1007), .ZN(n2537) );
  XNR2D1 U4081 ( .A1(s1_5_r[10]), .A2(W1_8_r[63]), .ZN(n2628) );
  AO21D1 U4082 ( .A1(n988), .A2(n2629), .B(n2628), .Z(
        dp_cluster_2_mult_485_C409_n296) );
  XNR2D1 U4083 ( .A1(n1010), .A2(n1371), .ZN(n2538) );
  XNR2D1 U4084 ( .A1(n1009), .A2(n1370), .ZN(n2627) );
  XNR2D1 U4085 ( .A1(n1009), .A2(n1372), .ZN(n2539) );
  XNR2D1 U4086 ( .A1(n1009), .A2(n1373), .ZN(n2540) );
  XNR2D1 U4087 ( .A1(n1009), .A2(n1374), .ZN(n2541) );
  XNR2D1 U4088 ( .A1(n1009), .A2(n1375), .ZN(n2542) );
  XNR2D1 U4089 ( .A1(n1009), .A2(n1376), .ZN(n2543) );
  XNR2D1 U4090 ( .A1(n1009), .A2(n1377), .ZN(n2544) );
  XNR2D1 U4091 ( .A1(n1009), .A2(n1378), .ZN(n2545) );
  XNR2D1 U4092 ( .A1(n1009), .A2(n1379), .ZN(n2546) );
  XNR2D1 U4093 ( .A1(n1009), .A2(n1380), .ZN(n2547) );
  XNR2D1 U4094 ( .A1(n1009), .A2(n1381), .ZN(n2548) );
  XNR2D1 U4095 ( .A1(n1009), .A2(n1382), .ZN(n2549) );
  XNR2D1 U4096 ( .A1(n1009), .A2(n1383), .ZN(n2550) );
  XNR2D1 U4097 ( .A1(n1091), .A2(n1010), .ZN(n2551) );
  XNR2D1 U4098 ( .A1(s1_5_r[8]), .A2(W1_8_r[63]), .ZN(n2552) );
  AO21D1 U4099 ( .A1(n986), .A2(n2569), .B(n2552), .Z(
        dp_cluster_2_mult_485_C409_n312) );
  XNR2D1 U4100 ( .A1(n1012), .A2(n1370), .ZN(n2553) );
  XNR2D1 U4101 ( .A1(n1012), .A2(n1371), .ZN(n2554) );
  XNR2D1 U4102 ( .A1(n1012), .A2(n1372), .ZN(n2555) );
  XNR2D1 U4103 ( .A1(n1012), .A2(n1373), .ZN(n2556) );
  XNR2D1 U4104 ( .A1(n1012), .A2(n1376), .ZN(n2559) );
  XNR2D1 U4105 ( .A1(n1012), .A2(n1377), .ZN(n2560) );
  XNR2D1 U4106 ( .A1(n1012), .A2(n1378), .ZN(n2561) );
  XNR2D1 U4107 ( .A1(n1012), .A2(n1379), .ZN(n2562) );
  XNR2D1 U4108 ( .A1(n1012), .A2(n1380), .ZN(n2563) );
  XNR2D1 U4109 ( .A1(n1012), .A2(n1381), .ZN(n2564) );
  XNR2D1 U4110 ( .A1(n1012), .A2(n1382), .ZN(n2565) );
  XNR2D1 U4111 ( .A1(n1012), .A2(n1383), .ZN(n2566) );
  XNR2D1 U4112 ( .A1(n1090), .A2(n1013), .ZN(n2568) );
  AO21D1 U4113 ( .A1(n984), .A2(n2587), .B(n2570), .Z(
        dp_cluster_2_mult_485_C409_n329) );
  XNR2D1 U4114 ( .A1(n1015), .A2(n1371), .ZN(n2572) );
  XNR2D1 U4115 ( .A1(n1015), .A2(n1372), .ZN(n2573) );
  XNR2D1 U4116 ( .A1(n1015), .A2(n1373), .ZN(n2574) );
  XNR2D1 U4117 ( .A1(n1015), .A2(n1374), .ZN(n2575) );
  XNR2D1 U4118 ( .A1(n1015), .A2(n1375), .ZN(n2576) );
  XNR2D1 U4119 ( .A1(n1015), .A2(n1376), .ZN(n2577) );
  XNR2D1 U4120 ( .A1(n1015), .A2(n1377), .ZN(n2578) );
  XNR2D1 U4121 ( .A1(n1015), .A2(n1378), .ZN(n2579) );
  XNR2D1 U4122 ( .A1(n1015), .A2(n1379), .ZN(n2580) );
  XNR2D1 U4123 ( .A1(n1015), .A2(n1380), .ZN(n2581) );
  XNR2D1 U4124 ( .A1(n1015), .A2(n1381), .ZN(n2582) );
  XNR2D1 U4125 ( .A1(n1015), .A2(n1382), .ZN(n2583) );
  XNR2D1 U4126 ( .A1(n1015), .A2(n1383), .ZN(n2584) );
  XNR2D1 U4127 ( .A1(n1090), .A2(n1016), .ZN(n2586) );
  AO21D1 U4128 ( .A1(n985), .A2(n2605), .B(n2588), .Z(
        dp_cluster_2_mult_485_C409_n345) );
  XNR2D1 U4129 ( .A1(n1018), .A2(n1371), .ZN(n2590) );
  XNR2D1 U4130 ( .A1(n1018), .A2(n1372), .ZN(n2591) );
  XNR2D1 U4131 ( .A1(n1018), .A2(n1373), .ZN(n2592) );
  XNR2D1 U4132 ( .A1(n1018), .A2(n1374), .ZN(n2593) );
  XNR2D1 U4133 ( .A1(n1018), .A2(n1375), .ZN(n2594) );
  XNR2D1 U4134 ( .A1(n1018), .A2(n1376), .ZN(n2595) );
  XNR2D1 U4135 ( .A1(n1018), .A2(n1377), .ZN(n2596) );
  XNR2D1 U4136 ( .A1(n1018), .A2(n1378), .ZN(n2597) );
  XNR2D1 U4137 ( .A1(n1018), .A2(n1379), .ZN(n2598) );
  XNR2D1 U4138 ( .A1(n1018), .A2(n1380), .ZN(n2599) );
  XNR2D1 U4139 ( .A1(n1018), .A2(n1381), .ZN(n2600) );
  XNR2D1 U4140 ( .A1(n1018), .A2(n1382), .ZN(n2601) );
  XNR2D1 U4141 ( .A1(n1018), .A2(n1383), .ZN(n2602) );
  XNR2D1 U4142 ( .A1(n1090), .A2(n1019), .ZN(n2604) );
  CKXOR2D1 U4143 ( .A1(n1112), .A2(W1_8_r[63]), .Z(n2606) );
  XNR2D1 U4144 ( .A1(n1112), .A2(W1_8_r[62]), .ZN(n2607) );
  MOAI22D1 U4145 ( .A1(n2607), .A2(n2621), .B1(n2606), .B2(s1_5_r[1]), .ZN(
        dp_cluster_2_mult_485_C409_n362) );
  XNR2D1 U4146 ( .A1(n1111), .A2(W1_8_r[61]), .ZN(n2608) );
  XNR2D1 U4147 ( .A1(n1112), .A2(W1_8_r[60]), .ZN(n2609) );
  XNR2D1 U4148 ( .A1(n1112), .A2(W1_8_r[59]), .ZN(n2610) );
  XNR2D1 U4149 ( .A1(n1111), .A2(W1_8_r[58]), .ZN(n2611) );
  XNR2D1 U4150 ( .A1(n1111), .A2(W1_8_r[57]), .ZN(n2612) );
  XNR2D1 U4151 ( .A1(n1111), .A2(W1_8_r[56]), .ZN(n2613) );
  XNR2D1 U4152 ( .A1(n1111), .A2(W1_8_r[55]), .ZN(n2614) );
  XNR2D1 U4153 ( .A1(n1111), .A2(W1_8_r[54]), .ZN(n2615) );
  XNR2D1 U4154 ( .A1(n1111), .A2(W1_8_r[53]), .ZN(n2616) );
  XNR2D1 U4155 ( .A1(n1111), .A2(W1_8_r[52]), .ZN(n2617) );
  XNR2D1 U4156 ( .A1(n1111), .A2(W1_8_r[51]), .ZN(n2618) );
  XNR2D1 U4157 ( .A1(n1111), .A2(W1_8_r[50]), .ZN(n2619) );
  XNR2D1 U4158 ( .A1(n1111), .A2(W1_8_r[49]), .ZN(n2620) );
  XNR2D1 U4159 ( .A1(W1_8_r[61]), .A2(s1_5_r[16]), .ZN(n2633) );
  XNR2D1 U4160 ( .A1(s1_5_r[14]), .A2(W1_8_r[63]), .ZN(n2634) );
  AN2XD1 U4161 ( .A1(n2642), .A2(n1135), .Z(n2641) );
  MAOI22D1 U4162 ( .A1(n2644), .A2(dp_cluster_2_N3), .B1(dp_cluster_2_N31), 
        .B2(n2643), .ZN(n2646) );
  AN2XD1 U4163 ( .A1(n2646), .A2(n1132), .Z(n2645) );
  MAOI22D1 U4164 ( .A1(n2648), .A2(dp_cluster_2_N5), .B1(dp_cluster_2_N33), 
        .B2(n2647), .ZN(n2650) );
  AN2XD1 U4165 ( .A1(n2650), .A2(n1128), .Z(n2649) );
  MAOI22D1 U4166 ( .A1(n2652), .A2(dp_cluster_2_N7), .B1(dp_cluster_2_N35), 
        .B2(n2651), .ZN(n2654) );
  AN2XD1 U4167 ( .A1(n2654), .A2(n1125), .Z(n2653) );
  MAOI22D1 U4168 ( .A1(n2656), .A2(dp_cluster_2_N9), .B1(dp_cluster_2_N37), 
        .B2(n2655), .ZN(n2658) );
  AN2XD1 U4169 ( .A1(n2658), .A2(n1121), .Z(n2657) );
  MAOI22D1 U4170 ( .A1(n2660), .A2(dp_cluster_2_N11), .B1(dp_cluster_2_N39), 
        .B2(n2659), .ZN(n2662) );
  AN2XD1 U4171 ( .A1(n2662), .A2(n1116), .Z(n2661) );
  XNR2D1 U4172 ( .A1(n1051), .A2(n1374), .ZN(n2701) );
  XNR2D1 U4173 ( .A1(n1051), .A2(s1_5_i[11]), .ZN(n2663) );
  XNR2D1 U4174 ( .A1(n1050), .A2(n1373), .ZN(n2700) );
  XNR2D1 U4175 ( .A1(s1_5_i[6]), .A2(W1_8_r[63]), .ZN(n2744) );
  XNR2D1 U4176 ( .A1(n1059), .A2(n1370), .ZN(n2745) );
  XNR2D1 U4177 ( .A1(n1059), .A2(s1_5_i[5]), .ZN(n2664) );
  XNR2D1 U4178 ( .A1(s1_5_i[4]), .A2(W1_8_r[63]), .ZN(n2762) );
  XNR2D1 U4179 ( .A1(n1062), .A2(n1370), .ZN(n2763) );
  XNR2D1 U4180 ( .A1(n1062), .A2(s1_5_i[3]), .ZN(n2665) );
  XNR2D1 U4181 ( .A1(n1056), .A2(n1375), .ZN(n2732) );
  XNR2D1 U4182 ( .A1(n1056), .A2(s1_5_i[7]), .ZN(n2666) );
  XNR2D1 U4183 ( .A1(n1056), .A2(n1374), .ZN(n2731) );
  XNR2D1 U4184 ( .A1(n1048), .A2(n1381), .ZN(n2694) );
  XNR2D1 U4185 ( .A1(n1048), .A2(s1_5_i[13]), .ZN(n2667) );
  XNR2D1 U4186 ( .A1(n1048), .A2(n1380), .ZN(n2693) );
  XNR2D1 U4187 ( .A1(n2669), .A2(n2668), .ZN(dp_cluster_3_mult_513_C415_n162)
         );
  XNR2D1 U4188 ( .A1(n1045), .A2(s1_5_i[15]), .ZN(n2670) );
  XNR2D1 U4189 ( .A1(n1053), .A2(s1_5_i[9]), .ZN(n2671) );
  XNR2D1 U4190 ( .A1(n1045), .A2(n1373), .ZN(n2672) );
  XNR2D1 U4191 ( .A1(s1_5_i[16]), .A2(W1_8_r[60]), .ZN(n2804) );
  XNR2D1 U4192 ( .A1(n1045), .A2(n1374), .ZN(n2673) );
  XNR2D1 U4193 ( .A1(n1045), .A2(n1375), .ZN(n2674) );
  XNR2D1 U4194 ( .A1(n1045), .A2(n1376), .ZN(n2675) );
  XNR2D1 U4195 ( .A1(n1045), .A2(n1377), .ZN(n2676) );
  XNR2D1 U4196 ( .A1(n1045), .A2(n1378), .ZN(n2677) );
  XNR2D1 U4197 ( .A1(n1045), .A2(n1379), .ZN(n2678) );
  XNR2D1 U4198 ( .A1(n1045), .A2(n1380), .ZN(n2679) );
  XNR2D1 U4199 ( .A1(n1045), .A2(n1381), .ZN(n2680) );
  XNR2D1 U4200 ( .A1(n1045), .A2(n1382), .ZN(n2681) );
  XNR2D1 U4201 ( .A1(n1045), .A2(n1383), .ZN(n2682) );
  XNR2D1 U4202 ( .A1(n1090), .A2(n1046), .ZN(n2683) );
  XNR2D1 U4203 ( .A1(n1047), .A2(n1371), .ZN(n2684) );
  XNR2D1 U4204 ( .A1(n1047), .A2(n1370), .ZN(n2811) );
  XNR2D1 U4205 ( .A1(n1047), .A2(n1372), .ZN(n2685) );
  XNR2D1 U4206 ( .A1(n1047), .A2(n1373), .ZN(n2686) );
  XNR2D1 U4207 ( .A1(n1048), .A2(n1374), .ZN(n2687) );
  XNR2D1 U4208 ( .A1(n1047), .A2(n1375), .ZN(n2688) );
  XNR2D1 U4209 ( .A1(n1047), .A2(n1376), .ZN(n2689) );
  XNR2D1 U4210 ( .A1(n1047), .A2(n1377), .ZN(n2690) );
  XNR2D1 U4211 ( .A1(n1047), .A2(n1378), .ZN(n2691) );
  XNR2D1 U4212 ( .A1(n1047), .A2(n1379), .ZN(n2692) );
  XNR2D1 U4213 ( .A1(n1047), .A2(n1382), .ZN(n2695) );
  XNR2D1 U4214 ( .A1(n1047), .A2(n1383), .ZN(n2696) );
  XNR2D1 U4215 ( .A1(n1089), .A2(n1049), .ZN(n2697) );
  XNR2D1 U4216 ( .A1(s1_5_i[12]), .A2(W1_8_r[63]), .ZN(n2798) );
  AO21D1 U4217 ( .A1(n989), .A2(n2799), .B(n2798), .Z(
        dp_cluster_3_mult_513_C415_n281) );
  XNR2D1 U4218 ( .A1(n1050), .A2(n1371), .ZN(n2698) );
  XNR2D1 U4219 ( .A1(n1050), .A2(n1370), .ZN(n2797) );
  XNR2D1 U4220 ( .A1(n1050), .A2(n1372), .ZN(n2699) );
  XNR2D1 U4221 ( .A1(n1050), .A2(n1375), .ZN(n2702) );
  XNR2D1 U4222 ( .A1(n1051), .A2(n1376), .ZN(n2703) );
  XNR2D1 U4223 ( .A1(n1050), .A2(n1377), .ZN(n2704) );
  XNR2D1 U4224 ( .A1(n1050), .A2(n1378), .ZN(n2705) );
  XNR2D1 U4225 ( .A1(n1050), .A2(n1379), .ZN(n2706) );
  XNR2D1 U4226 ( .A1(n1050), .A2(n1380), .ZN(n2707) );
  XNR2D1 U4227 ( .A1(n1050), .A2(n1381), .ZN(n2708) );
  XNR2D1 U4228 ( .A1(n1050), .A2(n1382), .ZN(n2709) );
  XNR2D1 U4229 ( .A1(n1050), .A2(n1383), .ZN(n2710) );
  XNR2D1 U4230 ( .A1(n1089), .A2(n1051), .ZN(n2711) );
  XNR2D1 U4231 ( .A1(s1_5_i[10]), .A2(W1_8_r[63]), .ZN(n2802) );
  AO21D1 U4232 ( .A1(n994), .A2(n2803), .B(n2802), .Z(
        dp_cluster_3_mult_513_C415_n296) );
  XNR2D1 U4233 ( .A1(n1053), .A2(n1371), .ZN(n2712) );
  XNR2D1 U4234 ( .A1(n1052), .A2(n1370), .ZN(n2801) );
  XNR2D1 U4235 ( .A1(n1052), .A2(n1372), .ZN(n2713) );
  XNR2D1 U4236 ( .A1(n1052), .A2(n1373), .ZN(n2714) );
  XNR2D1 U4237 ( .A1(n1052), .A2(n1374), .ZN(n2715) );
  XNR2D1 U4238 ( .A1(n1052), .A2(n1375), .ZN(n2716) );
  XNR2D1 U4239 ( .A1(n1053), .A2(n1376), .ZN(n2717) );
  XNR2D1 U4240 ( .A1(n1052), .A2(n1377), .ZN(n2718) );
  XNR2D1 U4241 ( .A1(n1052), .A2(n1378), .ZN(n2719) );
  XNR2D1 U4242 ( .A1(n1052), .A2(n1379), .ZN(n2720) );
  XNR2D1 U4243 ( .A1(n1052), .A2(n1380), .ZN(n2721) );
  XNR2D1 U4244 ( .A1(n1052), .A2(n1381), .ZN(n2722) );
  XNR2D1 U4245 ( .A1(n1052), .A2(n1382), .ZN(n2723) );
  XNR2D1 U4246 ( .A1(n1052), .A2(n1383), .ZN(n2724) );
  XNR2D1 U4247 ( .A1(n1089), .A2(n1054), .ZN(n2725) );
  XNR2D1 U4248 ( .A1(s1_5_i[8]), .A2(W1_8_r[63]), .ZN(n2726) );
  AO21D1 U4249 ( .A1(n992), .A2(n2743), .B(n2726), .Z(
        dp_cluster_3_mult_513_C415_n312) );
  XNR2D1 U4250 ( .A1(n1055), .A2(n1370), .ZN(n2727) );
  XNR2D1 U4251 ( .A1(n1055), .A2(n1371), .ZN(n2728) );
  XNR2D1 U4252 ( .A1(n1055), .A2(n1372), .ZN(n2729) );
  XNR2D1 U4253 ( .A1(n1055), .A2(n1373), .ZN(n2730) );
  XNR2D1 U4254 ( .A1(n1056), .A2(n1376), .ZN(n2733) );
  XNR2D1 U4255 ( .A1(n1055), .A2(n1377), .ZN(n2734) );
  XNR2D1 U4256 ( .A1(n1055), .A2(n1378), .ZN(n2735) );
  XNR2D1 U4257 ( .A1(n1055), .A2(n1379), .ZN(n2736) );
  XNR2D1 U4258 ( .A1(n1055), .A2(n1380), .ZN(n2737) );
  XNR2D1 U4259 ( .A1(n1055), .A2(n1381), .ZN(n2738) );
  XNR2D1 U4260 ( .A1(n1055), .A2(n1382), .ZN(n2739) );
  XNR2D1 U4261 ( .A1(n1055), .A2(n1383), .ZN(n2740) );
  XNR2D1 U4262 ( .A1(n1089), .A2(n1057), .ZN(n2742) );
  AO21D1 U4263 ( .A1(n990), .A2(n2761), .B(n2744), .Z(
        dp_cluster_3_mult_513_C415_n329) );
  XNR2D1 U4264 ( .A1(n1058), .A2(n1371), .ZN(n2746) );
  XNR2D1 U4265 ( .A1(n1058), .A2(n1372), .ZN(n2747) );
  XNR2D1 U4266 ( .A1(n1058), .A2(n1373), .ZN(n2748) );
  XNR2D1 U4267 ( .A1(n1058), .A2(n1374), .ZN(n2749) );
  XNR2D1 U4268 ( .A1(n1058), .A2(n1375), .ZN(n2750) );
  XNR2D1 U4269 ( .A1(n1059), .A2(n1376), .ZN(n2751) );
  XNR2D1 U4270 ( .A1(n1058), .A2(n1377), .ZN(n2752) );
  XNR2D1 U4271 ( .A1(n1058), .A2(n1378), .ZN(n2753) );
  XNR2D1 U4272 ( .A1(n1058), .A2(n1379), .ZN(n2754) );
  XNR2D1 U4273 ( .A1(n1058), .A2(n1380), .ZN(n2755) );
  XNR2D1 U4274 ( .A1(n1058), .A2(n1381), .ZN(n2756) );
  XNR2D1 U4275 ( .A1(n1058), .A2(n1382), .ZN(n2757) );
  XNR2D1 U4276 ( .A1(n1058), .A2(n1383), .ZN(n2758) );
  XNR2D1 U4277 ( .A1(n1089), .A2(n1060), .ZN(n2760) );
  AO21D1 U4278 ( .A1(n991), .A2(n2779), .B(n2762), .Z(
        dp_cluster_3_mult_513_C415_n345) );
  XNR2D1 U4279 ( .A1(n1061), .A2(n1371), .ZN(n2764) );
  XNR2D1 U4280 ( .A1(n1061), .A2(n1372), .ZN(n2765) );
  XNR2D1 U4281 ( .A1(n1061), .A2(n1373), .ZN(n2766) );
  XNR2D1 U4282 ( .A1(n1061), .A2(n1374), .ZN(n2767) );
  XNR2D1 U4283 ( .A1(n1061), .A2(n1375), .ZN(n2768) );
  XNR2D1 U4284 ( .A1(n1062), .A2(n1376), .ZN(n2769) );
  XNR2D1 U4285 ( .A1(n1061), .A2(n1377), .ZN(n2770) );
  XNR2D1 U4286 ( .A1(n1061), .A2(n1378), .ZN(n2771) );
  XNR2D1 U4287 ( .A1(n1061), .A2(n1379), .ZN(n2772) );
  XNR2D1 U4288 ( .A1(n1061), .A2(n1380), .ZN(n2773) );
  XNR2D1 U4289 ( .A1(n1061), .A2(n1381), .ZN(n2774) );
  XNR2D1 U4290 ( .A1(n1061), .A2(n1382), .ZN(n2775) );
  XNR2D1 U4291 ( .A1(n1061), .A2(n1383), .ZN(n2776) );
  XNR2D1 U4292 ( .A1(n1089), .A2(n1063), .ZN(n2778) );
  CKXOR2D1 U4293 ( .A1(n1105), .A2(W1_8_r[63]), .Z(n2780) );
  XNR2D1 U4294 ( .A1(n1105), .A2(W1_8_r[62]), .ZN(n2781) );
  MOAI22D1 U4295 ( .A1(n2781), .A2(n2795), .B1(n2780), .B2(s1_5_i[1]), .ZN(
        dp_cluster_3_mult_513_C415_n362) );
  XNR2D1 U4296 ( .A1(n1104), .A2(W1_8_r[61]), .ZN(n2782) );
  XNR2D1 U4297 ( .A1(n1104), .A2(W1_8_r[60]), .ZN(n2783) );
  XNR2D1 U4298 ( .A1(n1104), .A2(W1_8_r[59]), .ZN(n2784) );
  XNR2D1 U4299 ( .A1(n1104), .A2(W1_8_r[58]), .ZN(n2785) );
  XNR2D1 U4300 ( .A1(n1104), .A2(W1_8_r[57]), .ZN(n2786) );
  XNR2D1 U4301 ( .A1(n1104), .A2(W1_8_r[56]), .ZN(n2787) );
  XNR2D1 U4302 ( .A1(n1104), .A2(W1_8_r[55]), .ZN(n2788) );
  XNR2D1 U4303 ( .A1(n1104), .A2(W1_8_r[54]), .ZN(n2789) );
  XNR2D1 U4304 ( .A1(n1104), .A2(W1_8_r[53]), .ZN(n2790) );
  XNR2D1 U4305 ( .A1(n1104), .A2(W1_8_r[52]), .ZN(n2791) );
  XNR2D1 U4306 ( .A1(n1104), .A2(W1_8_r[51]), .ZN(n2792) );
  XNR2D1 U4307 ( .A1(n1104), .A2(W1_8_r[50]), .ZN(n2793) );
  XNR2D1 U4308 ( .A1(n1105), .A2(W1_8_r[49]), .ZN(n2794) );
  XNR2D1 U4309 ( .A1(W1_8_r[61]), .A2(s1_5_i[16]), .ZN(n2807) );
  XNR2D1 U4310 ( .A1(s1_5_i[14]), .A2(W1_8_r[63]), .ZN(n2808) );
  XNR2D1 U4311 ( .A1(n1007), .A2(n1404), .ZN(n2853) );
  XNR2D1 U4312 ( .A1(n1007), .A2(s1_5_r[11]), .ZN(n2815) );
  XNR2D1 U4313 ( .A1(n1006), .A2(n1403), .ZN(n2852) );
  XNR2D1 U4314 ( .A1(s1_5_r[6]), .A2(W1_8_i[63]), .ZN(n2896) );
  XNR2D1 U4315 ( .A1(n1015), .A2(n1400), .ZN(n2897) );
  XNR2D1 U4316 ( .A1(n1015), .A2(s1_5_r[5]), .ZN(n2816) );
  XNR2D1 U4317 ( .A1(s1_5_r[4]), .A2(W1_8_i[63]), .ZN(n2914) );
  XNR2D1 U4318 ( .A1(n1018), .A2(n1400), .ZN(n2915) );
  XNR2D1 U4319 ( .A1(n1018), .A2(s1_5_r[3]), .ZN(n2817) );
  XNR2D1 U4320 ( .A1(n1012), .A2(n1405), .ZN(n2884) );
  XNR2D1 U4321 ( .A1(n1012), .A2(s1_5_r[7]), .ZN(n2818) );
  XNR2D1 U4322 ( .A1(n1012), .A2(n1404), .ZN(n2883) );
  XNR2D1 U4323 ( .A1(n1004), .A2(n1411), .ZN(n2846) );
  XNR2D1 U4324 ( .A1(n1004), .A2(s1_5_r[13]), .ZN(n2819) );
  XNR2D1 U4325 ( .A1(n1004), .A2(n1410), .ZN(n2845) );
  XNR2D1 U4326 ( .A1(n2821), .A2(n2820), .ZN(dp_cluster_3_mult_512_C415_n162)
         );
  XNR2D1 U4327 ( .A1(n1001), .A2(s1_5_r[15]), .ZN(n2822) );
  XNR2D1 U4328 ( .A1(n1009), .A2(s1_5_r[9]), .ZN(n2823) );
  XNR2D1 U4329 ( .A1(n1001), .A2(n1403), .ZN(n2824) );
  XNR2D1 U4330 ( .A1(s1_5_r[16]), .A2(W1_8_i[60]), .ZN(n2956) );
  XNR2D1 U4331 ( .A1(n1001), .A2(n1404), .ZN(n2825) );
  XNR2D1 U4332 ( .A1(n1001), .A2(n1405), .ZN(n2826) );
  XNR2D1 U4333 ( .A1(n1001), .A2(n1406), .ZN(n2827) );
  XNR2D1 U4334 ( .A1(n1001), .A2(n1407), .ZN(n2828) );
  XNR2D1 U4335 ( .A1(n1001), .A2(n1408), .ZN(n2829) );
  XNR2D1 U4336 ( .A1(n1001), .A2(n1409), .ZN(n2830) );
  XNR2D1 U4337 ( .A1(n1001), .A2(n1410), .ZN(n2831) );
  XNR2D1 U4338 ( .A1(n1001), .A2(n1411), .ZN(n2832) );
  XNR2D1 U4339 ( .A1(n1001), .A2(n1412), .ZN(n2833) );
  XNR2D1 U4340 ( .A1(n1001), .A2(n1413), .ZN(n2834) );
  XNR2D1 U4341 ( .A1(n1096), .A2(n1002), .ZN(n2835) );
  XNR2D1 U4342 ( .A1(n1003), .A2(n1401), .ZN(n2836) );
  XNR2D1 U4343 ( .A1(n1003), .A2(n1400), .ZN(n2963) );
  XNR2D1 U4344 ( .A1(n1003), .A2(n1402), .ZN(n2837) );
  XNR2D1 U4345 ( .A1(n1003), .A2(n1403), .ZN(n2838) );
  XNR2D1 U4346 ( .A1(n1004), .A2(n1404), .ZN(n2839) );
  XNR2D1 U4347 ( .A1(n1003), .A2(n1405), .ZN(n2840) );
  XNR2D1 U4348 ( .A1(n1003), .A2(n1406), .ZN(n2841) );
  XNR2D1 U4349 ( .A1(n1003), .A2(n1407), .ZN(n2842) );
  XNR2D1 U4350 ( .A1(n1003), .A2(n1408), .ZN(n2843) );
  XNR2D1 U4351 ( .A1(n1003), .A2(n1409), .ZN(n2844) );
  XNR2D1 U4352 ( .A1(n1003), .A2(n1412), .ZN(n2847) );
  XNR2D1 U4353 ( .A1(n1003), .A2(n1413), .ZN(n2848) );
  XNR2D1 U4354 ( .A1(n1095), .A2(n1005), .ZN(n2849) );
  XNR2D1 U4355 ( .A1(s1_5_r[12]), .A2(W1_8_i[63]), .ZN(n2950) );
  AO21D1 U4356 ( .A1(n995), .A2(n2951), .B(n2950), .Z(
        dp_cluster_3_mult_512_C415_n281) );
  XNR2D1 U4357 ( .A1(n1006), .A2(n1401), .ZN(n2850) );
  XNR2D1 U4358 ( .A1(n1006), .A2(n1400), .ZN(n2949) );
  XNR2D1 U4359 ( .A1(n1006), .A2(n1402), .ZN(n2851) );
  XNR2D1 U4360 ( .A1(n1006), .A2(n1405), .ZN(n2854) );
  XNR2D1 U4361 ( .A1(n1007), .A2(n1406), .ZN(n2855) );
  XNR2D1 U4362 ( .A1(n1006), .A2(n1407), .ZN(n2856) );
  XNR2D1 U4363 ( .A1(n1006), .A2(n1408), .ZN(n2857) );
  XNR2D1 U4364 ( .A1(n1006), .A2(n1409), .ZN(n2858) );
  XNR2D1 U4365 ( .A1(n1006), .A2(n1410), .ZN(n2859) );
  XNR2D1 U4366 ( .A1(n1006), .A2(n1411), .ZN(n2860) );
  XNR2D1 U4367 ( .A1(n1006), .A2(n1412), .ZN(n2861) );
  XNR2D1 U4368 ( .A1(n1006), .A2(n1413), .ZN(n2862) );
  XNR2D1 U4369 ( .A1(n1095), .A2(n1007), .ZN(n2863) );
  XNR2D1 U4370 ( .A1(s1_5_r[10]), .A2(W1_8_i[63]), .ZN(n2954) );
  AO21D1 U4371 ( .A1(n1000), .A2(n2955), .B(n2954), .Z(
        dp_cluster_3_mult_512_C415_n296) );
  XNR2D1 U4372 ( .A1(n1009), .A2(n1401), .ZN(n2864) );
  XNR2D1 U4373 ( .A1(n1008), .A2(n1400), .ZN(n2953) );
  XNR2D1 U4374 ( .A1(n1008), .A2(n1402), .ZN(n2865) );
  XNR2D1 U4375 ( .A1(n1008), .A2(n1403), .ZN(n2866) );
  XNR2D1 U4376 ( .A1(n1008), .A2(n1404), .ZN(n2867) );
  XNR2D1 U4377 ( .A1(n1008), .A2(n1405), .ZN(n2868) );
  XNR2D1 U4378 ( .A1(n1009), .A2(n1406), .ZN(n2869) );
  XNR2D1 U4379 ( .A1(n1008), .A2(n1407), .ZN(n2870) );
  XNR2D1 U4380 ( .A1(n1008), .A2(n1408), .ZN(n2871) );
  XNR2D1 U4381 ( .A1(n1008), .A2(n1409), .ZN(n2872) );
  XNR2D1 U4382 ( .A1(n1008), .A2(n1410), .ZN(n2873) );
  XNR2D1 U4383 ( .A1(n1008), .A2(n1411), .ZN(n2874) );
  XNR2D1 U4384 ( .A1(n1008), .A2(n1412), .ZN(n2875) );
  XNR2D1 U4385 ( .A1(n1008), .A2(n1413), .ZN(n2876) );
  XNR2D1 U4386 ( .A1(n1095), .A2(n1010), .ZN(n2877) );
  XNR2D1 U4387 ( .A1(s1_5_r[8]), .A2(W1_8_i[63]), .ZN(n2878) );
  AO21D1 U4388 ( .A1(n998), .A2(n2895), .B(n2878), .Z(
        dp_cluster_3_mult_512_C415_n312) );
  XNR2D1 U4389 ( .A1(n1011), .A2(n1400), .ZN(n2879) );
  XNR2D1 U4390 ( .A1(n1011), .A2(n1401), .ZN(n2880) );
  XNR2D1 U4391 ( .A1(n1011), .A2(n1402), .ZN(n2881) );
  XNR2D1 U4392 ( .A1(n1011), .A2(n1403), .ZN(n2882) );
  XNR2D1 U4393 ( .A1(n1012), .A2(n1406), .ZN(n2885) );
  XNR2D1 U4394 ( .A1(n1011), .A2(n1407), .ZN(n2886) );
  XNR2D1 U4395 ( .A1(n1011), .A2(n1408), .ZN(n2887) );
  XNR2D1 U4396 ( .A1(n1011), .A2(n1409), .ZN(n2888) );
  XNR2D1 U4397 ( .A1(n1011), .A2(n1410), .ZN(n2889) );
  XNR2D1 U4398 ( .A1(n1011), .A2(n1411), .ZN(n2890) );
  XNR2D1 U4399 ( .A1(n1011), .A2(n1412), .ZN(n2891) );
  XNR2D1 U4400 ( .A1(n1011), .A2(n1413), .ZN(n2892) );
  XNR2D1 U4401 ( .A1(n1095), .A2(n1013), .ZN(n2894) );
  AO21D1 U4402 ( .A1(n996), .A2(n2913), .B(n2896), .Z(
        dp_cluster_3_mult_512_C415_n329) );
  XNR2D1 U4403 ( .A1(n1014), .A2(n1401), .ZN(n2898) );
  XNR2D1 U4404 ( .A1(n1014), .A2(n1402), .ZN(n2899) );
  XNR2D1 U4405 ( .A1(n1014), .A2(n1403), .ZN(n2900) );
  XNR2D1 U4406 ( .A1(n1014), .A2(n1404), .ZN(n2901) );
  XNR2D1 U4407 ( .A1(n1014), .A2(n1405), .ZN(n2902) );
  XNR2D1 U4408 ( .A1(n1015), .A2(n1406), .ZN(n2903) );
  XNR2D1 U4409 ( .A1(n1014), .A2(n1407), .ZN(n2904) );
  XNR2D1 U4410 ( .A1(n1014), .A2(n1408), .ZN(n2905) );
  XNR2D1 U4411 ( .A1(n1014), .A2(n1409), .ZN(n2906) );
  XNR2D1 U4412 ( .A1(n1014), .A2(n1410), .ZN(n2907) );
  XNR2D1 U4413 ( .A1(n1014), .A2(n1411), .ZN(n2908) );
  XNR2D1 U4414 ( .A1(n1014), .A2(n1412), .ZN(n2909) );
  XNR2D1 U4415 ( .A1(n1014), .A2(n1413), .ZN(n2910) );
  XNR2D1 U4416 ( .A1(n1095), .A2(n1016), .ZN(n2912) );
  AO21D1 U4417 ( .A1(n997), .A2(n2931), .B(n2914), .Z(
        dp_cluster_3_mult_512_C415_n345) );
  XNR2D1 U4418 ( .A1(n1017), .A2(n1401), .ZN(n2916) );
  XNR2D1 U4419 ( .A1(n1017), .A2(n1402), .ZN(n2917) );
  XNR2D1 U4420 ( .A1(n1017), .A2(n1403), .ZN(n2918) );
  XNR2D1 U4421 ( .A1(n1017), .A2(n1404), .ZN(n2919) );
  XNR2D1 U4422 ( .A1(n1017), .A2(n1405), .ZN(n2920) );
  XNR2D1 U4423 ( .A1(n1018), .A2(n1406), .ZN(n2921) );
  XNR2D1 U4424 ( .A1(n1017), .A2(n1407), .ZN(n2922) );
  XNR2D1 U4425 ( .A1(n1017), .A2(n1408), .ZN(n2923) );
  XNR2D1 U4426 ( .A1(n1017), .A2(n1409), .ZN(n2924) );
  XNR2D1 U4427 ( .A1(n1017), .A2(n1410), .ZN(n2925) );
  XNR2D1 U4428 ( .A1(n1017), .A2(n1411), .ZN(n2926) );
  XNR2D1 U4429 ( .A1(n1017), .A2(n1412), .ZN(n2927) );
  XNR2D1 U4430 ( .A1(n1017), .A2(n1413), .ZN(n2928) );
  XNR2D1 U4431 ( .A1(n1095), .A2(n1019), .ZN(n2930) );
  CKXOR2D1 U4432 ( .A1(n1111), .A2(W1_8_i[63]), .Z(n2932) );
  XNR2D1 U4433 ( .A1(n1111), .A2(W1_8_i[62]), .ZN(n2933) );
  MOAI22D1 U4434 ( .A1(n2933), .A2(n2947), .B1(n2932), .B2(s1_5_r[1]), .ZN(
        dp_cluster_3_mult_512_C415_n362) );
  XNR2D1 U4435 ( .A1(n1110), .A2(W1_8_i[61]), .ZN(n2934) );
  XNR2D1 U4436 ( .A1(n1110), .A2(W1_8_i[60]), .ZN(n2935) );
  XNR2D1 U4437 ( .A1(n1110), .A2(W1_8_i[59]), .ZN(n2936) );
  XNR2D1 U4438 ( .A1(n1110), .A2(W1_8_i[58]), .ZN(n2937) );
  XNR2D1 U4439 ( .A1(n1110), .A2(W1_8_i[57]), .ZN(n2938) );
  XNR2D1 U4440 ( .A1(n1110), .A2(W1_8_i[56]), .ZN(n2939) );
  XNR2D1 U4441 ( .A1(n1110), .A2(W1_8_i[55]), .ZN(n2940) );
  XNR2D1 U4442 ( .A1(n1110), .A2(W1_8_i[54]), .ZN(n2941) );
  XNR2D1 U4443 ( .A1(n1110), .A2(W1_8_i[53]), .ZN(n2942) );
  XNR2D1 U4444 ( .A1(n1110), .A2(W1_8_i[52]), .ZN(n2943) );
  XNR2D1 U4445 ( .A1(n1110), .A2(W1_8_i[51]), .ZN(n2944) );
  XNR2D1 U4446 ( .A1(n1110), .A2(W1_8_i[50]), .ZN(n2945) );
  XNR2D1 U4447 ( .A1(n1111), .A2(W1_8_i[49]), .ZN(n2946) );
  XNR2D1 U4448 ( .A1(W1_8_i[61]), .A2(s1_5_r[16]), .ZN(n2959) );
  XNR2D1 U4449 ( .A1(s1_5_r[14]), .A2(W1_8_i[63]), .ZN(n2960) );
endmodule

