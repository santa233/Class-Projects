
module alu2_tj ( a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p );
  input a, b, c, d, e, f, g, h, i, j;
  output k, l, m, n, o, p;
  wire   n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712;

  IV U369 ( .A(g), .Z(n608) );
  IV U370 ( .A(a), .Z(n581) );
  AN2 U371 ( .A(n608), .B(n581), .Z(n398) );
  IV U372 ( .A(h), .Z(n637) );
  OR2 U373 ( .A(j), .B(n637), .Z(n459) );
  AN2 U374 ( .A(e), .B(f), .Z(n692) );
  IV U375 ( .A(n692), .Z(n537) );
  OR2 U376 ( .A(n537), .B(h), .Z(n364) );
  AN2 U377 ( .A(n459), .B(n364), .Z(n365) );
  OR2 U378 ( .A(n365), .B(n608), .Z(n367) );
  OR2 U379 ( .A(n608), .B(h), .Z(n504) );
  IV U380 ( .A(n504), .Z(n385) );
  IV U381 ( .A(e), .Z(n659) );
  AN2 U382 ( .A(n659), .B(f), .Z(n662) );
  IV U383 ( .A(n662), .Z(n625) );
  OR2 U384 ( .A(n385), .B(n625), .Z(n366) );
  AN2 U385 ( .A(n367), .B(n366), .Z(n479) );
  OR2 U386 ( .A(c), .B(n479), .Z(n371) );
  IV U387 ( .A(j), .Z(n376) );
  OR2 U388 ( .A(n376), .B(g), .Z(n413) );
  IV U389 ( .A(n413), .Z(n497) );
  IV U390 ( .A(f), .Z(n630) );
  AN2 U391 ( .A(n630), .B(e), .Z(n689) );
  AN2 U392 ( .A(n459), .B(n689), .Z(n368) );
  IV U393 ( .A(n368), .Z(n369) );
  OR2 U394 ( .A(n497), .B(n369), .Z(n490) );
  IV U395 ( .A(c), .Z(n446) );
  AN2 U396 ( .A(n581), .B(n446), .Z(n706) );
  OR2 U397 ( .A(n490), .B(n706), .Z(n370) );
  AN2 U398 ( .A(n371), .B(n370), .Z(n375) );
  AN2 U399 ( .A(j), .B(h), .Z(n536) );
  AN2 U400 ( .A(n608), .B(n536), .Z(n690) );
  IV U401 ( .A(n690), .Z(n503) );
  AN2 U402 ( .A(n659), .B(n630), .Z(n564) );
  IV U403 ( .A(n564), .Z(n513) );
  OR2 U404 ( .A(n513), .B(n504), .Z(n372) );
  AN2 U405 ( .A(n503), .B(n372), .Z(n373) );
  OR2 U406 ( .A(n581), .B(n446), .Z(n468) );
  OR2 U407 ( .A(n373), .B(n468), .Z(n374) );
  AN2 U408 ( .A(n375), .B(n374), .Z(n418) );
  IV U409 ( .A(n398), .Z(n377) );
  AN2 U410 ( .A(n377), .B(n376), .Z(n383) );
  OR2 U411 ( .A(c), .B(n581), .Z(n449) );
  OR2 U412 ( .A(n446), .B(a), .Z(n499) );
  OR2 U413 ( .A(n504), .B(n499), .Z(n378) );
  AN2 U414 ( .A(n449), .B(n378), .Z(n379) );
  OR2 U415 ( .A(n379), .B(n630), .Z(n380) );
  AN2 U416 ( .A(j), .B(n380), .Z(n381) );
  OR2 U417 ( .A(n381), .B(e), .Z(n382) );
  OR2 U418 ( .A(n383), .B(n382), .Z(n384) );
  AN2 U419 ( .A(n418), .B(n384), .Z(n576) );
  IV U420 ( .A(n576), .Z(n575) );
  IV U421 ( .A(n468), .Z(n707) );
  AN2 U422 ( .A(n608), .B(n707), .Z(n552) );
  AN2 U423 ( .A(j), .B(n385), .Z(n590) );
  AN2 U424 ( .A(n575), .B(a), .Z(n681) );
  AN2 U425 ( .A(n692), .B(n681), .Z(n426) );
  AN2 U426 ( .A(n707), .B(n689), .Z(n387) );
  AN2 U427 ( .A(n576), .B(n564), .Z(n386) );
  OR2 U428 ( .A(n387), .B(n386), .Z(n388) );
  OR2 U429 ( .A(n426), .B(n388), .Z(n389) );
  AN2 U430 ( .A(n590), .B(n389), .Z(n391) );
  AN2 U431 ( .A(n662), .B(n536), .Z(n518) );
  AN2 U432 ( .A(n518), .B(n575), .Z(n390) );
  OR2 U433 ( .A(n391), .B(n390), .Z(n551) );
  IV U434 ( .A(n551), .Z(n589) );
  AN2 U435 ( .A(n689), .B(n589), .Z(n392) );
  OR2 U436 ( .A(n552), .B(n392), .Z(n549) );
  OR2 U437 ( .A(n575), .B(n549), .Z(n393) );
  IV U438 ( .A(n393), .Z(n395) );
  AN2 U439 ( .A(n575), .B(n549), .Z(n523) );
  OR2 U440 ( .A(n523), .B(f), .Z(n394) );
  OR2 U441 ( .A(n395), .B(n394), .Z(n396) );
  AN2 U442 ( .A(g), .B(n396), .Z(n397) );
  OR2 U443 ( .A(n398), .B(n397), .Z(n401) );
  AN2 U444 ( .A(n551), .B(a), .Z(n657) );
  AN2 U445 ( .A(n589), .B(n537), .Z(n399) );
  OR2 U446 ( .A(n657), .B(n399), .Z(n400) );
  AN2 U447 ( .A(n401), .B(n400), .Z(n404) );
  AN2 U448 ( .A(g), .B(n576), .Z(n660) );
  IV U449 ( .A(n660), .Z(n546) );
  OR2 U450 ( .A(g), .B(n576), .Z(n402) );
  AN2 U451 ( .A(n546), .B(n402), .Z(n440) );
  OR2 U452 ( .A(n625), .B(n440), .Z(n403) );
  AN2 U453 ( .A(n404), .B(n403), .Z(n406) );
  AN2 U454 ( .A(n637), .B(j), .Z(n672) );
  IV U455 ( .A(n672), .Z(n405) );
  OR2 U456 ( .A(n406), .B(n405), .Z(n417) );
  OR2 U457 ( .A(n692), .B(n575), .Z(n407) );
  AN2 U458 ( .A(a), .B(n407), .Z(n411) );
  AN2 U459 ( .A(g), .B(n536), .Z(n582) );
  OR2 U460 ( .A(a), .B(n407), .Z(n408) );
  AN2 U461 ( .A(n582), .B(n408), .Z(n409) );
  IV U462 ( .A(n409), .Z(n410) );
  OR2 U463 ( .A(n411), .B(n410), .Z(n415) );
  IV U464 ( .A(n689), .Z(n622) );
  OR2 U465 ( .A(n499), .B(n622), .Z(n445) );
  AN2 U466 ( .A(n445), .B(n449), .Z(n412) );
  OR2 U467 ( .A(n413), .B(n412), .Z(n414) );
  AN2 U468 ( .A(n415), .B(n414), .Z(n416) );
  AN2 U469 ( .A(n417), .B(n416), .Z(n424) );
  OR2 U470 ( .A(n707), .B(n589), .Z(n421) );
  AN2 U471 ( .A(n692), .B(n418), .Z(n419) );
  IV U472 ( .A(n419), .Z(n420) );
  AN2 U473 ( .A(n421), .B(n420), .Z(n422) );
  OR2 U474 ( .A(n503), .B(n422), .Z(n423) );
  AN2 U475 ( .A(n424), .B(n423), .Z(n600) );
  IV U476 ( .A(i), .Z(n462) );
  AN2 U477 ( .A(j), .B(n462), .Z(n425) );
  AN2 U478 ( .A(n600), .B(n425), .Z(n467) );
  IV U479 ( .A(n426), .Z(n437) );
  OR2 U480 ( .A(n625), .B(a), .Z(n427) );
  AN2 U481 ( .A(n622), .B(n427), .Z(n428) );
  OR2 U482 ( .A(n428), .B(n504), .Z(n429) );
  AN2 U483 ( .A(n429), .B(n446), .Z(n432) );
  OR2 U484 ( .A(e), .B(g), .Z(n483) );
  OR2 U485 ( .A(n483), .B(n576), .Z(n430) );
  AN2 U486 ( .A(c), .B(n430), .Z(n431) );
  OR2 U487 ( .A(n432), .B(n431), .Z(n435) );
  OR2 U488 ( .A(n608), .B(n625), .Z(n433) );
  OR2 U489 ( .A(n468), .B(n433), .Z(n434) );
  AN2 U490 ( .A(n435), .B(n434), .Z(n436) );
  AN2 U491 ( .A(n437), .B(n436), .Z(n439) );
  OR2 U492 ( .A(h), .B(n622), .Z(n610) );
  OR2 U493 ( .A(n610), .B(n575), .Z(n438) );
  AN2 U494 ( .A(n439), .B(n438), .Z(n442) );
  OR2 U495 ( .A(n513), .B(n440), .Z(n441) );
  AN2 U496 ( .A(n442), .B(n441), .Z(n443) );
  OR2 U497 ( .A(n443), .B(j), .Z(n458) );
  AN2 U498 ( .A(n608), .B(n672), .Z(n530) );
  AN2 U499 ( .A(n692), .B(n530), .Z(n444) );
  IV U500 ( .A(n444), .Z(n642) );
  OR2 U501 ( .A(n445), .B(g), .Z(n448) );
  OR2 U502 ( .A(n625), .B(n446), .Z(n447) );
  AN2 U503 ( .A(n448), .B(n447), .Z(n454) );
  AN2 U504 ( .A(n468), .B(f), .Z(n452) );
  AN2 U505 ( .A(n576), .B(n449), .Z(n450) );
  AN2 U506 ( .A(n450), .B(n630), .Z(n451) );
  OR2 U507 ( .A(n452), .B(n451), .Z(n453) );
  AN2 U508 ( .A(n454), .B(n453), .Z(n455) );
  OR2 U509 ( .A(n459), .B(n455), .Z(n456) );
  AN2 U510 ( .A(n642), .B(n456), .Z(n457) );
  AN2 U511 ( .A(n458), .B(n457), .Z(n461) );
  AN2 U512 ( .A(n608), .B(n513), .Z(n534) );
  OR2 U513 ( .A(n534), .B(n459), .Z(n643) );
  OR2 U514 ( .A(n581), .B(n643), .Z(n460) );
  AN2 U515 ( .A(n461), .B(n460), .Z(n464) );
  OR2 U516 ( .A(n600), .B(n462), .Z(n463) );
  AN2 U517 ( .A(n464), .B(n463), .Z(n465) );
  IV U518 ( .A(n465), .Z(n466) );
  OR2 U519 ( .A(n467), .B(n466), .Z(k) );
  IV U520 ( .A(b), .Z(n644) );
  IV U521 ( .A(d), .Z(n626) );
  OR2 U522 ( .A(n644), .B(n626), .Z(n628) );
  IV U523 ( .A(n628), .Z(n709) );
  OR2 U524 ( .A(n709), .B(n468), .Z(n469) );
  AN2 U525 ( .A(n497), .B(n469), .Z(n472) );
  OR2 U526 ( .A(b), .B(n626), .Z(n493) );
  OR2 U527 ( .A(d), .B(n644), .Z(n629) );
  AN2 U528 ( .A(n493), .B(n629), .Z(n710) );
  IV U529 ( .A(n710), .Z(n470) );
  AN2 U530 ( .A(n472), .B(n470), .Z(n475) );
  OR2 U531 ( .A(b), .B(d), .Z(n686) );
  IV U532 ( .A(n686), .Z(n489) );
  AN2 U533 ( .A(n690), .B(n489), .Z(n471) );
  OR2 U534 ( .A(n472), .B(n471), .Z(n473) );
  AN2 U535 ( .A(n707), .B(n473), .Z(n474) );
  OR2 U536 ( .A(n475), .B(n474), .Z(n529) );
  AN2 U537 ( .A(n629), .B(n499), .Z(n478) );
  IV U538 ( .A(n499), .Z(n495) );
  AN2 U539 ( .A(n495), .B(n686), .Z(n476) );
  OR2 U540 ( .A(n476), .B(n625), .Z(n477) );
  OR2 U541 ( .A(n478), .B(n477), .Z(n488) );
  OR2 U542 ( .A(d), .B(n479), .Z(n482) );
  AN2 U543 ( .A(a), .B(n582), .Z(n580) );
  AN2 U544 ( .A(n580), .B(n564), .Z(n480) );
  IV U545 ( .A(n480), .Z(n481) );
  AN2 U546 ( .A(n482), .B(n481), .Z(n486) );
  OR2 U547 ( .A(n483), .B(j), .Z(n484) );
  OR2 U548 ( .A(b), .B(n484), .Z(n485) );
  AN2 U549 ( .A(n486), .B(n485), .Z(n487) );
  AN2 U550 ( .A(n488), .B(n487), .Z(n492) );
  OR2 U551 ( .A(n490), .B(n489), .Z(n491) );
  AN2 U552 ( .A(n492), .B(n491), .Z(n512) );
  IV U553 ( .A(n590), .Z(n498) );
  OR2 U554 ( .A(n493), .B(n625), .Z(n494) );
  OR2 U555 ( .A(n495), .B(n494), .Z(n496) );
  OR2 U556 ( .A(n498), .B(n496), .Z(n510) );
  AN2 U557 ( .A(n692), .B(n497), .Z(n678) );
  IV U558 ( .A(n678), .Z(n502) );
  OR2 U559 ( .A(n499), .B(n498), .Z(n500) );
  OR2 U560 ( .A(e), .B(n500), .Z(n501) );
  AN2 U561 ( .A(n502), .B(n501), .Z(n507) );
  AN2 U562 ( .A(n504), .B(n503), .Z(n505) );
  OR2 U563 ( .A(n513), .B(n505), .Z(n506) );
  AN2 U564 ( .A(n507), .B(n506), .Z(n508) );
  OR2 U565 ( .A(n628), .B(n508), .Z(n509) );
  AN2 U566 ( .A(n510), .B(n509), .Z(n511) );
  AN2 U567 ( .A(n512), .B(n511), .Z(n661) );
  IV U568 ( .A(n661), .Z(n613) );
  OR2 U569 ( .A(g), .B(n628), .Z(n652) );
  AN2 U570 ( .A(n689), .B(n709), .Z(n516) );
  OR2 U571 ( .A(n513), .B(n613), .Z(n602) );
  IV U572 ( .A(n602), .Z(n514) );
  AN2 U573 ( .A(n613), .B(b), .Z(n683) );
  AN2 U574 ( .A(n692), .B(n683), .Z(n619) );
  OR2 U575 ( .A(n514), .B(n619), .Z(n515) );
  OR2 U576 ( .A(n516), .B(n515), .Z(n517) );
  AN2 U577 ( .A(n590), .B(n517), .Z(n520) );
  OR2 U578 ( .A(b), .B(n613), .Z(n680) );
  AN2 U579 ( .A(n518), .B(n680), .Z(n519) );
  OR2 U580 ( .A(n520), .B(n519), .Z(n655) );
  OR2 U581 ( .A(n655), .B(n622), .Z(n521) );
  AN2 U582 ( .A(n652), .B(n521), .Z(n553) );
  IV U583 ( .A(n553), .Z(n522) );
  AN2 U584 ( .A(n613), .B(n522), .Z(n524) );
  OR2 U585 ( .A(n523), .B(n524), .Z(n669) );
  IV U586 ( .A(n669), .Z(n526) );
  AN2 U587 ( .A(n524), .B(n523), .Z(n525) );
  OR2 U588 ( .A(n526), .B(n525), .Z(n527) );
  AN2 U589 ( .A(n590), .B(n527), .Z(n528) );
  OR2 U590 ( .A(n529), .B(n528), .Z(n532) );
  AN2 U591 ( .A(d), .B(n530), .Z(n531) );
  OR2 U592 ( .A(n532), .B(n531), .Z(n533) );
  AN2 U593 ( .A(n689), .B(n533), .Z(n599) );
  IV U594 ( .A(n655), .Z(n653) );
  OR2 U595 ( .A(n653), .B(n657), .Z(n565) );
  IV U596 ( .A(n565), .Z(n544) );
  IV U597 ( .A(n534), .Z(n535) );
  AN2 U598 ( .A(n536), .B(n535), .Z(n538) );
  AN2 U599 ( .A(n538), .B(n537), .Z(n685) );
  IV U600 ( .A(n681), .Z(n539) );
  AN2 U601 ( .A(n539), .B(n661), .Z(n541) );
  AN2 U602 ( .A(n681), .B(n613), .Z(n540) );
  OR2 U603 ( .A(n541), .B(n540), .Z(n571) );
  IV U604 ( .A(n571), .Z(n542) );
  AN2 U605 ( .A(n685), .B(n542), .Z(n543) );
  OR2 U606 ( .A(n544), .B(n543), .Z(n545) );
  AN2 U607 ( .A(n644), .B(n545), .Z(n563) );
  AN2 U608 ( .A(n672), .B(n546), .Z(n547) );
  AN2 U609 ( .A(n613), .B(n547), .Z(n558) );
  AN2 U610 ( .A(n652), .B(n655), .Z(n548) );
  OR2 U611 ( .A(n549), .B(n548), .Z(n550) );
  AN2 U612 ( .A(n690), .B(n550), .Z(n556) );
  AN2 U613 ( .A(n551), .B(n655), .Z(n584) );
  AN2 U614 ( .A(n552), .B(n584), .Z(n705) );
  AN2 U615 ( .A(n553), .B(n705), .Z(n554) );
  IV U616 ( .A(n554), .Z(n555) );
  AN2 U617 ( .A(n556), .B(n555), .Z(n557) );
  OR2 U618 ( .A(n558), .B(n557), .Z(n560) );
  AN2 U619 ( .A(n661), .B(n576), .Z(n679) );
  AN2 U620 ( .A(n590), .B(n679), .Z(n559) );
  OR2 U621 ( .A(n560), .B(n559), .Z(n561) );
  AN2 U622 ( .A(n662), .B(n561), .Z(n562) );
  OR2 U623 ( .A(n563), .B(n562), .Z(n597) );
  AN2 U624 ( .A(n565), .B(n564), .Z(n568) );
  AN2 U625 ( .A(n657), .B(n653), .Z(n566) );
  IV U626 ( .A(n566), .Z(n567) );
  AN2 U627 ( .A(n568), .B(n567), .Z(n569) );
  OR2 U628 ( .A(n569), .B(n608), .Z(n570) );
  AN2 U629 ( .A(n672), .B(n570), .Z(n573) );
  AN2 U630 ( .A(n571), .B(n685), .Z(n572) );
  OR2 U631 ( .A(n573), .B(n572), .Z(n574) );
  AN2 U632 ( .A(b), .B(n574), .Z(n595) );
  OR2 U633 ( .A(n661), .B(n575), .Z(n578) );
  OR2 U634 ( .A(n576), .B(n613), .Z(n577) );
  AN2 U635 ( .A(n578), .B(n577), .Z(n579) );
  AN2 U636 ( .A(n690), .B(n579), .Z(n588) );
  AN2 U637 ( .A(n580), .B(b), .Z(n586) );
  AN2 U638 ( .A(n582), .B(n581), .Z(n583) );
  AN2 U639 ( .A(n583), .B(n644), .Z(n693) );
  OR2 U640 ( .A(n693), .B(n584), .Z(n585) );
  OR2 U641 ( .A(n586), .B(n585), .Z(n587) );
  OR2 U642 ( .A(n588), .B(n587), .Z(n592) );
  AN2 U643 ( .A(n589), .B(n653), .Z(n664) );
  AN2 U644 ( .A(n590), .B(n664), .Z(n591) );
  OR2 U645 ( .A(n592), .B(n591), .Z(n593) );
  AN2 U646 ( .A(n692), .B(n593), .Z(n594) );
  OR2 U647 ( .A(n595), .B(n594), .Z(n596) );
  OR2 U648 ( .A(n597), .B(n596), .Z(n598) );
  OR2 U649 ( .A(n599), .B(n598), .Z(n674) );
  OR2 U650 ( .A(i), .B(n600), .Z(n673) );
  AN2 U651 ( .A(n674), .B(n673), .Z(n651) );
  OR2 U652 ( .A(n625), .B(n628), .Z(n601) );
  AN2 U653 ( .A(n602), .B(n601), .Z(n607) );
  OR2 U654 ( .A(n625), .B(b), .Z(n603) );
  AN2 U655 ( .A(n622), .B(n603), .Z(n604) );
  OR2 U656 ( .A(n604), .B(d), .Z(n605) );
  OR2 U657 ( .A(h), .B(n605), .Z(n606) );
  AN2 U658 ( .A(n607), .B(n606), .Z(n609) );
  OR2 U659 ( .A(n609), .B(n608), .Z(n618) );
  AN2 U660 ( .A(n661), .B(n610), .Z(n616) );
  AN2 U661 ( .A(n626), .B(f), .Z(n611) );
  OR2 U662 ( .A(e), .B(n611), .Z(n612) );
  AN2 U663 ( .A(n613), .B(n612), .Z(n614) );
  OR2 U664 ( .A(n614), .B(g), .Z(n615) );
  OR2 U665 ( .A(n616), .B(n615), .Z(n617) );
  AN2 U666 ( .A(n618), .B(n617), .Z(n621) );
  IV U667 ( .A(n619), .Z(n620) );
  AN2 U668 ( .A(n621), .B(n620), .Z(n639) );
  OR2 U669 ( .A(g), .B(n622), .Z(n623) );
  OR2 U670 ( .A(n623), .B(b), .Z(n624) );
  AN2 U671 ( .A(n625), .B(n624), .Z(n627) );
  OR2 U672 ( .A(n627), .B(n626), .Z(n635) );
  AN2 U673 ( .A(n628), .B(f), .Z(n633) );
  AN2 U674 ( .A(n661), .B(n629), .Z(n631) );
  AN2 U675 ( .A(n631), .B(n630), .Z(n632) );
  OR2 U676 ( .A(n633), .B(n632), .Z(n634) );
  AN2 U677 ( .A(n635), .B(n634), .Z(n636) );
  OR2 U678 ( .A(n637), .B(n636), .Z(n638) );
  AN2 U679 ( .A(n639), .B(n638), .Z(n640) );
  OR2 U680 ( .A(n640), .B(j), .Z(n641) );
  AN2 U681 ( .A(n642), .B(n641), .Z(n646) );
  OR2 U682 ( .A(n644), .B(n643), .Z(n645) );
  AN2 U683 ( .A(n646), .B(n645), .Z(n648) );
  OR2 U684 ( .A(n674), .B(n673), .Z(n647) );
  AN2 U685 ( .A(n648), .B(n647), .Z(n649) );
  IV U686 ( .A(n649), .Z(n650) );
  OR2 U687 ( .A(n651), .B(n650), .Z(l) );
  OR2 U688 ( .A(n653), .B(n652), .Z(n654) );
  IV U689 ( .A(n654), .Z(n703) );
  AN2 U690 ( .A(b), .B(n655), .Z(n656) );
  OR2 U691 ( .A(n657), .B(n656), .Z(n658) );
  AN2 U692 ( .A(n659), .B(n658), .Z(n668) );
  AN2 U693 ( .A(n661), .B(n660), .Z(n663) );
  AN2 U694 ( .A(n663), .B(n662), .Z(n666) );
  AN2 U695 ( .A(n664), .B(n692), .Z(n665) );
  OR2 U696 ( .A(n666), .B(n665), .Z(n667) );
  OR2 U697 ( .A(n668), .B(n667), .Z(n670) );
  OR2 U698 ( .A(n670), .B(n669), .Z(n671) );
  AN2 U699 ( .A(n672), .B(n671), .Z(n677) );
  IV U700 ( .A(n673), .Z(n675) );
  AN2 U701 ( .A(n675), .B(n674), .Z(n676) );
  OR2 U702 ( .A(n677), .B(n676), .Z(n701) );
  AN2 U703 ( .A(n679), .B(n678), .Z(n699) );
  AN2 U704 ( .A(n681), .B(n680), .Z(n682) );
  OR2 U705 ( .A(n683), .B(n682), .Z(n684) );
  AN2 U706 ( .A(n685), .B(n684), .Z(n697) );
  AN2 U707 ( .A(n707), .B(n686), .Z(n687) );
  OR2 U708 ( .A(n709), .B(n687), .Z(n688) );
  AN2 U709 ( .A(n689), .B(n688), .Z(n691) );
  AN2 U710 ( .A(n691), .B(n690), .Z(n695) );
  AN2 U711 ( .A(n693), .B(n692), .Z(n694) );
  OR2 U712 ( .A(n695), .B(n694), .Z(n696) );
  OR2 U713 ( .A(n697), .B(n696), .Z(n698) );
  OR2 U714 ( .A(n699), .B(n698), .Z(n700) );
  OR2 U715 ( .A(n701), .B(n700), .Z(n702) );
  OR2 U716 ( .A(n703), .B(n702), .Z(n704) );
  OR2 U717 ( .A(n705), .B(n704), .Z(o) );
  OR2 U718 ( .A(n707), .B(n706), .Z(n708) );
  AN2 U719 ( .A(n710), .B(n708), .Z(p) );
  IV U720 ( .A(n709), .Z(n711) );
  IV U721 ( .A(n711), .Z(n) );
  IV U722 ( .A(n710), .Z(n712) );
  IV U723 ( .A(n712), .Z(m) );
  
  
endmodule

